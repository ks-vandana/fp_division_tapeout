magic
tech sky130A
magscale 1 2
timestamp 1700930463
<< obsli1 >>
rect 1104 2159 158884 157777
<< obsm1 >>
rect 1104 2128 159054 157888
<< metal2 >>
rect 2686 159200 2742 160000
rect 7102 159200 7158 160000
rect 11518 159200 11574 160000
rect 15934 159200 15990 160000
rect 20350 159200 20406 160000
rect 24766 159200 24822 160000
rect 29182 159200 29238 160000
rect 33598 159200 33654 160000
rect 38014 159200 38070 160000
rect 42430 159200 42486 160000
rect 46846 159200 46902 160000
rect 51262 159200 51318 160000
rect 55678 159200 55734 160000
rect 60094 159200 60150 160000
rect 64510 159200 64566 160000
rect 68926 159200 68982 160000
rect 73342 159200 73398 160000
rect 77758 159200 77814 160000
rect 82174 159200 82230 160000
rect 86590 159200 86646 160000
rect 91006 159200 91062 160000
rect 95422 159200 95478 160000
rect 99838 159200 99894 160000
rect 104254 159200 104310 160000
rect 108670 159200 108726 160000
rect 113086 159200 113142 160000
rect 117502 159200 117558 160000
rect 121918 159200 121974 160000
rect 126334 159200 126390 160000
rect 130750 159200 130806 160000
rect 135166 159200 135222 160000
rect 139582 159200 139638 160000
rect 143998 159200 144054 160000
rect 148414 159200 148470 160000
rect 152830 159200 152886 160000
rect 157246 159200 157302 160000
rect 11886 0 11942 800
rect 12162 0 12218 800
rect 12438 0 12494 800
rect 12714 0 12770 800
rect 12990 0 13046 800
rect 13266 0 13322 800
rect 13542 0 13598 800
rect 13818 0 13874 800
rect 14094 0 14150 800
rect 14370 0 14426 800
rect 14646 0 14702 800
rect 14922 0 14978 800
rect 15198 0 15254 800
rect 15474 0 15530 800
rect 15750 0 15806 800
rect 16026 0 16082 800
rect 16302 0 16358 800
rect 16578 0 16634 800
rect 16854 0 16910 800
rect 17130 0 17186 800
rect 17406 0 17462 800
rect 17682 0 17738 800
rect 17958 0 18014 800
rect 18234 0 18290 800
rect 18510 0 18566 800
rect 18786 0 18842 800
rect 19062 0 19118 800
rect 19338 0 19394 800
rect 19614 0 19670 800
rect 19890 0 19946 800
rect 20166 0 20222 800
rect 20442 0 20498 800
rect 20718 0 20774 800
rect 20994 0 21050 800
rect 21270 0 21326 800
rect 21546 0 21602 800
rect 21822 0 21878 800
rect 22098 0 22154 800
rect 22374 0 22430 800
rect 22650 0 22706 800
rect 22926 0 22982 800
rect 23202 0 23258 800
rect 23478 0 23534 800
rect 23754 0 23810 800
rect 24030 0 24086 800
rect 24306 0 24362 800
rect 24582 0 24638 800
rect 24858 0 24914 800
rect 25134 0 25190 800
rect 25410 0 25466 800
rect 25686 0 25742 800
rect 25962 0 26018 800
rect 26238 0 26294 800
rect 26514 0 26570 800
rect 26790 0 26846 800
rect 27066 0 27122 800
rect 27342 0 27398 800
rect 27618 0 27674 800
rect 27894 0 27950 800
rect 28170 0 28226 800
rect 28446 0 28502 800
rect 28722 0 28778 800
rect 28998 0 29054 800
rect 29274 0 29330 800
rect 29550 0 29606 800
rect 29826 0 29882 800
rect 30102 0 30158 800
rect 30378 0 30434 800
rect 30654 0 30710 800
rect 30930 0 30986 800
rect 31206 0 31262 800
rect 31482 0 31538 800
rect 31758 0 31814 800
rect 32034 0 32090 800
rect 32310 0 32366 800
rect 32586 0 32642 800
rect 32862 0 32918 800
rect 33138 0 33194 800
rect 33414 0 33470 800
rect 33690 0 33746 800
rect 33966 0 34022 800
rect 34242 0 34298 800
rect 34518 0 34574 800
rect 34794 0 34850 800
rect 35070 0 35126 800
rect 35346 0 35402 800
rect 35622 0 35678 800
rect 35898 0 35954 800
rect 36174 0 36230 800
rect 36450 0 36506 800
rect 36726 0 36782 800
rect 37002 0 37058 800
rect 37278 0 37334 800
rect 37554 0 37610 800
rect 37830 0 37886 800
rect 38106 0 38162 800
rect 38382 0 38438 800
rect 38658 0 38714 800
rect 38934 0 38990 800
rect 39210 0 39266 800
rect 39486 0 39542 800
rect 39762 0 39818 800
rect 40038 0 40094 800
rect 40314 0 40370 800
rect 40590 0 40646 800
rect 40866 0 40922 800
rect 41142 0 41198 800
rect 41418 0 41474 800
rect 41694 0 41750 800
rect 41970 0 42026 800
rect 42246 0 42302 800
rect 42522 0 42578 800
rect 42798 0 42854 800
rect 43074 0 43130 800
rect 43350 0 43406 800
rect 43626 0 43682 800
rect 43902 0 43958 800
rect 44178 0 44234 800
rect 44454 0 44510 800
rect 44730 0 44786 800
rect 45006 0 45062 800
rect 45282 0 45338 800
rect 45558 0 45614 800
rect 45834 0 45890 800
rect 46110 0 46166 800
rect 46386 0 46442 800
rect 46662 0 46718 800
rect 46938 0 46994 800
rect 47214 0 47270 800
rect 47490 0 47546 800
rect 47766 0 47822 800
rect 48042 0 48098 800
rect 48318 0 48374 800
rect 48594 0 48650 800
rect 48870 0 48926 800
rect 49146 0 49202 800
rect 49422 0 49478 800
rect 49698 0 49754 800
rect 49974 0 50030 800
rect 50250 0 50306 800
rect 50526 0 50582 800
rect 50802 0 50858 800
rect 51078 0 51134 800
rect 51354 0 51410 800
rect 51630 0 51686 800
rect 51906 0 51962 800
rect 52182 0 52238 800
rect 52458 0 52514 800
rect 52734 0 52790 800
rect 53010 0 53066 800
rect 53286 0 53342 800
rect 53562 0 53618 800
rect 53838 0 53894 800
rect 54114 0 54170 800
rect 54390 0 54446 800
rect 54666 0 54722 800
rect 54942 0 54998 800
rect 55218 0 55274 800
rect 55494 0 55550 800
rect 55770 0 55826 800
rect 56046 0 56102 800
rect 56322 0 56378 800
rect 56598 0 56654 800
rect 56874 0 56930 800
rect 57150 0 57206 800
rect 57426 0 57482 800
rect 57702 0 57758 800
rect 57978 0 58034 800
rect 58254 0 58310 800
rect 58530 0 58586 800
rect 58806 0 58862 800
rect 59082 0 59138 800
rect 59358 0 59414 800
rect 59634 0 59690 800
rect 59910 0 59966 800
rect 60186 0 60242 800
rect 60462 0 60518 800
rect 60738 0 60794 800
rect 61014 0 61070 800
rect 61290 0 61346 800
rect 61566 0 61622 800
rect 61842 0 61898 800
rect 62118 0 62174 800
rect 62394 0 62450 800
rect 62670 0 62726 800
rect 62946 0 63002 800
rect 63222 0 63278 800
rect 63498 0 63554 800
rect 63774 0 63830 800
rect 64050 0 64106 800
rect 64326 0 64382 800
rect 64602 0 64658 800
rect 64878 0 64934 800
rect 65154 0 65210 800
rect 65430 0 65486 800
rect 65706 0 65762 800
rect 65982 0 66038 800
rect 66258 0 66314 800
rect 66534 0 66590 800
rect 66810 0 66866 800
rect 67086 0 67142 800
rect 67362 0 67418 800
rect 67638 0 67694 800
rect 67914 0 67970 800
rect 68190 0 68246 800
rect 68466 0 68522 800
rect 68742 0 68798 800
rect 69018 0 69074 800
rect 69294 0 69350 800
rect 69570 0 69626 800
rect 69846 0 69902 800
rect 70122 0 70178 800
rect 70398 0 70454 800
rect 70674 0 70730 800
rect 70950 0 71006 800
rect 71226 0 71282 800
rect 71502 0 71558 800
rect 71778 0 71834 800
rect 72054 0 72110 800
rect 72330 0 72386 800
rect 72606 0 72662 800
rect 72882 0 72938 800
rect 73158 0 73214 800
rect 73434 0 73490 800
rect 73710 0 73766 800
rect 73986 0 74042 800
rect 74262 0 74318 800
rect 74538 0 74594 800
rect 74814 0 74870 800
rect 75090 0 75146 800
rect 75366 0 75422 800
rect 75642 0 75698 800
rect 75918 0 75974 800
rect 76194 0 76250 800
rect 76470 0 76526 800
rect 76746 0 76802 800
rect 77022 0 77078 800
rect 77298 0 77354 800
rect 77574 0 77630 800
rect 77850 0 77906 800
rect 78126 0 78182 800
rect 78402 0 78458 800
rect 78678 0 78734 800
rect 78954 0 79010 800
rect 79230 0 79286 800
rect 79506 0 79562 800
rect 79782 0 79838 800
rect 80058 0 80114 800
rect 80334 0 80390 800
rect 80610 0 80666 800
rect 80886 0 80942 800
rect 81162 0 81218 800
rect 81438 0 81494 800
rect 81714 0 81770 800
rect 81990 0 82046 800
rect 82266 0 82322 800
rect 82542 0 82598 800
rect 82818 0 82874 800
rect 83094 0 83150 800
rect 83370 0 83426 800
rect 83646 0 83702 800
rect 83922 0 83978 800
rect 84198 0 84254 800
rect 84474 0 84530 800
rect 84750 0 84806 800
rect 85026 0 85082 800
rect 85302 0 85358 800
rect 85578 0 85634 800
rect 85854 0 85910 800
rect 86130 0 86186 800
rect 86406 0 86462 800
rect 86682 0 86738 800
rect 86958 0 87014 800
rect 87234 0 87290 800
rect 87510 0 87566 800
rect 87786 0 87842 800
rect 88062 0 88118 800
rect 88338 0 88394 800
rect 88614 0 88670 800
rect 88890 0 88946 800
rect 89166 0 89222 800
rect 89442 0 89498 800
rect 89718 0 89774 800
rect 89994 0 90050 800
rect 90270 0 90326 800
rect 90546 0 90602 800
rect 90822 0 90878 800
rect 91098 0 91154 800
rect 91374 0 91430 800
rect 91650 0 91706 800
rect 91926 0 91982 800
rect 92202 0 92258 800
rect 92478 0 92534 800
rect 92754 0 92810 800
rect 93030 0 93086 800
rect 93306 0 93362 800
rect 93582 0 93638 800
rect 93858 0 93914 800
rect 94134 0 94190 800
rect 94410 0 94466 800
rect 94686 0 94742 800
rect 94962 0 95018 800
rect 95238 0 95294 800
rect 95514 0 95570 800
rect 95790 0 95846 800
rect 96066 0 96122 800
rect 96342 0 96398 800
rect 96618 0 96674 800
rect 96894 0 96950 800
rect 97170 0 97226 800
rect 97446 0 97502 800
rect 97722 0 97778 800
rect 97998 0 98054 800
rect 98274 0 98330 800
rect 98550 0 98606 800
rect 98826 0 98882 800
rect 99102 0 99158 800
rect 99378 0 99434 800
rect 99654 0 99710 800
rect 99930 0 99986 800
rect 100206 0 100262 800
rect 100482 0 100538 800
rect 100758 0 100814 800
rect 101034 0 101090 800
rect 101310 0 101366 800
rect 101586 0 101642 800
rect 101862 0 101918 800
rect 102138 0 102194 800
rect 102414 0 102470 800
rect 102690 0 102746 800
rect 102966 0 103022 800
rect 103242 0 103298 800
rect 103518 0 103574 800
rect 103794 0 103850 800
rect 104070 0 104126 800
rect 104346 0 104402 800
rect 104622 0 104678 800
rect 104898 0 104954 800
rect 105174 0 105230 800
rect 105450 0 105506 800
rect 105726 0 105782 800
rect 106002 0 106058 800
rect 106278 0 106334 800
rect 106554 0 106610 800
rect 106830 0 106886 800
rect 107106 0 107162 800
rect 107382 0 107438 800
rect 107658 0 107714 800
rect 107934 0 107990 800
rect 108210 0 108266 800
rect 108486 0 108542 800
rect 108762 0 108818 800
rect 109038 0 109094 800
rect 109314 0 109370 800
rect 109590 0 109646 800
rect 109866 0 109922 800
rect 110142 0 110198 800
rect 110418 0 110474 800
rect 110694 0 110750 800
rect 110970 0 111026 800
rect 111246 0 111302 800
rect 111522 0 111578 800
rect 111798 0 111854 800
rect 112074 0 112130 800
rect 112350 0 112406 800
rect 112626 0 112682 800
rect 112902 0 112958 800
rect 113178 0 113234 800
rect 113454 0 113510 800
rect 113730 0 113786 800
rect 114006 0 114062 800
rect 114282 0 114338 800
rect 114558 0 114614 800
rect 114834 0 114890 800
rect 115110 0 115166 800
rect 115386 0 115442 800
rect 115662 0 115718 800
rect 115938 0 115994 800
rect 116214 0 116270 800
rect 116490 0 116546 800
rect 116766 0 116822 800
rect 117042 0 117098 800
rect 117318 0 117374 800
rect 117594 0 117650 800
rect 117870 0 117926 800
rect 118146 0 118202 800
rect 118422 0 118478 800
rect 118698 0 118754 800
rect 118974 0 119030 800
rect 119250 0 119306 800
rect 119526 0 119582 800
rect 119802 0 119858 800
rect 120078 0 120134 800
rect 120354 0 120410 800
rect 120630 0 120686 800
rect 120906 0 120962 800
rect 121182 0 121238 800
rect 121458 0 121514 800
rect 121734 0 121790 800
rect 122010 0 122066 800
rect 122286 0 122342 800
rect 122562 0 122618 800
rect 122838 0 122894 800
rect 123114 0 123170 800
rect 123390 0 123446 800
rect 123666 0 123722 800
rect 123942 0 123998 800
rect 124218 0 124274 800
rect 124494 0 124550 800
rect 124770 0 124826 800
rect 125046 0 125102 800
rect 125322 0 125378 800
rect 125598 0 125654 800
rect 125874 0 125930 800
rect 126150 0 126206 800
rect 126426 0 126482 800
rect 126702 0 126758 800
rect 126978 0 127034 800
rect 127254 0 127310 800
rect 127530 0 127586 800
rect 127806 0 127862 800
rect 128082 0 128138 800
rect 128358 0 128414 800
rect 128634 0 128690 800
rect 128910 0 128966 800
rect 129186 0 129242 800
rect 129462 0 129518 800
rect 129738 0 129794 800
rect 130014 0 130070 800
rect 130290 0 130346 800
rect 130566 0 130622 800
rect 130842 0 130898 800
rect 131118 0 131174 800
rect 131394 0 131450 800
rect 131670 0 131726 800
rect 131946 0 132002 800
rect 132222 0 132278 800
rect 132498 0 132554 800
rect 132774 0 132830 800
rect 133050 0 133106 800
rect 133326 0 133382 800
rect 133602 0 133658 800
rect 133878 0 133934 800
rect 134154 0 134210 800
rect 134430 0 134486 800
rect 134706 0 134762 800
rect 134982 0 135038 800
rect 135258 0 135314 800
rect 135534 0 135590 800
rect 135810 0 135866 800
rect 136086 0 136142 800
rect 136362 0 136418 800
rect 136638 0 136694 800
rect 136914 0 136970 800
rect 137190 0 137246 800
rect 137466 0 137522 800
rect 137742 0 137798 800
rect 138018 0 138074 800
rect 138294 0 138350 800
rect 138570 0 138626 800
rect 138846 0 138902 800
rect 139122 0 139178 800
rect 139398 0 139454 800
rect 139674 0 139730 800
rect 139950 0 140006 800
rect 140226 0 140282 800
rect 140502 0 140558 800
rect 140778 0 140834 800
rect 141054 0 141110 800
rect 141330 0 141386 800
rect 141606 0 141662 800
rect 141882 0 141938 800
rect 142158 0 142214 800
rect 142434 0 142490 800
rect 142710 0 142766 800
rect 142986 0 143042 800
rect 143262 0 143318 800
rect 143538 0 143594 800
rect 143814 0 143870 800
rect 144090 0 144146 800
rect 144366 0 144422 800
rect 144642 0 144698 800
rect 144918 0 144974 800
rect 145194 0 145250 800
rect 145470 0 145526 800
rect 145746 0 145802 800
rect 146022 0 146078 800
rect 146298 0 146354 800
rect 146574 0 146630 800
rect 146850 0 146906 800
rect 147126 0 147182 800
rect 147402 0 147458 800
rect 147678 0 147734 800
rect 147954 0 148010 800
<< obsm2 >>
rect 1492 159144 2630 159338
rect 2798 159144 7046 159338
rect 7214 159144 11462 159338
rect 11630 159144 15878 159338
rect 16046 159144 20294 159338
rect 20462 159144 24710 159338
rect 24878 159144 29126 159338
rect 29294 159144 33542 159338
rect 33710 159144 37958 159338
rect 38126 159144 42374 159338
rect 42542 159144 46790 159338
rect 46958 159144 51206 159338
rect 51374 159144 55622 159338
rect 55790 159144 60038 159338
rect 60206 159144 64454 159338
rect 64622 159144 68870 159338
rect 69038 159144 73286 159338
rect 73454 159144 77702 159338
rect 77870 159144 82118 159338
rect 82286 159144 86534 159338
rect 86702 159144 90950 159338
rect 91118 159144 95366 159338
rect 95534 159144 99782 159338
rect 99950 159144 104198 159338
rect 104366 159144 108614 159338
rect 108782 159144 113030 159338
rect 113198 159144 117446 159338
rect 117614 159144 121862 159338
rect 122030 159144 126278 159338
rect 126446 159144 130694 159338
rect 130862 159144 135110 159338
rect 135278 159144 139526 159338
rect 139694 159144 143942 159338
rect 144110 159144 148358 159338
rect 148526 159144 152774 159338
rect 152942 159144 157190 159338
rect 157358 159144 159050 159338
rect 1492 856 159050 159144
rect 1492 800 11830 856
rect 11998 800 12106 856
rect 12274 800 12382 856
rect 12550 800 12658 856
rect 12826 800 12934 856
rect 13102 800 13210 856
rect 13378 800 13486 856
rect 13654 800 13762 856
rect 13930 800 14038 856
rect 14206 800 14314 856
rect 14482 800 14590 856
rect 14758 800 14866 856
rect 15034 800 15142 856
rect 15310 800 15418 856
rect 15586 800 15694 856
rect 15862 800 15970 856
rect 16138 800 16246 856
rect 16414 800 16522 856
rect 16690 800 16798 856
rect 16966 800 17074 856
rect 17242 800 17350 856
rect 17518 800 17626 856
rect 17794 800 17902 856
rect 18070 800 18178 856
rect 18346 800 18454 856
rect 18622 800 18730 856
rect 18898 800 19006 856
rect 19174 800 19282 856
rect 19450 800 19558 856
rect 19726 800 19834 856
rect 20002 800 20110 856
rect 20278 800 20386 856
rect 20554 800 20662 856
rect 20830 800 20938 856
rect 21106 800 21214 856
rect 21382 800 21490 856
rect 21658 800 21766 856
rect 21934 800 22042 856
rect 22210 800 22318 856
rect 22486 800 22594 856
rect 22762 800 22870 856
rect 23038 800 23146 856
rect 23314 800 23422 856
rect 23590 800 23698 856
rect 23866 800 23974 856
rect 24142 800 24250 856
rect 24418 800 24526 856
rect 24694 800 24802 856
rect 24970 800 25078 856
rect 25246 800 25354 856
rect 25522 800 25630 856
rect 25798 800 25906 856
rect 26074 800 26182 856
rect 26350 800 26458 856
rect 26626 800 26734 856
rect 26902 800 27010 856
rect 27178 800 27286 856
rect 27454 800 27562 856
rect 27730 800 27838 856
rect 28006 800 28114 856
rect 28282 800 28390 856
rect 28558 800 28666 856
rect 28834 800 28942 856
rect 29110 800 29218 856
rect 29386 800 29494 856
rect 29662 800 29770 856
rect 29938 800 30046 856
rect 30214 800 30322 856
rect 30490 800 30598 856
rect 30766 800 30874 856
rect 31042 800 31150 856
rect 31318 800 31426 856
rect 31594 800 31702 856
rect 31870 800 31978 856
rect 32146 800 32254 856
rect 32422 800 32530 856
rect 32698 800 32806 856
rect 32974 800 33082 856
rect 33250 800 33358 856
rect 33526 800 33634 856
rect 33802 800 33910 856
rect 34078 800 34186 856
rect 34354 800 34462 856
rect 34630 800 34738 856
rect 34906 800 35014 856
rect 35182 800 35290 856
rect 35458 800 35566 856
rect 35734 800 35842 856
rect 36010 800 36118 856
rect 36286 800 36394 856
rect 36562 800 36670 856
rect 36838 800 36946 856
rect 37114 800 37222 856
rect 37390 800 37498 856
rect 37666 800 37774 856
rect 37942 800 38050 856
rect 38218 800 38326 856
rect 38494 800 38602 856
rect 38770 800 38878 856
rect 39046 800 39154 856
rect 39322 800 39430 856
rect 39598 800 39706 856
rect 39874 800 39982 856
rect 40150 800 40258 856
rect 40426 800 40534 856
rect 40702 800 40810 856
rect 40978 800 41086 856
rect 41254 800 41362 856
rect 41530 800 41638 856
rect 41806 800 41914 856
rect 42082 800 42190 856
rect 42358 800 42466 856
rect 42634 800 42742 856
rect 42910 800 43018 856
rect 43186 800 43294 856
rect 43462 800 43570 856
rect 43738 800 43846 856
rect 44014 800 44122 856
rect 44290 800 44398 856
rect 44566 800 44674 856
rect 44842 800 44950 856
rect 45118 800 45226 856
rect 45394 800 45502 856
rect 45670 800 45778 856
rect 45946 800 46054 856
rect 46222 800 46330 856
rect 46498 800 46606 856
rect 46774 800 46882 856
rect 47050 800 47158 856
rect 47326 800 47434 856
rect 47602 800 47710 856
rect 47878 800 47986 856
rect 48154 800 48262 856
rect 48430 800 48538 856
rect 48706 800 48814 856
rect 48982 800 49090 856
rect 49258 800 49366 856
rect 49534 800 49642 856
rect 49810 800 49918 856
rect 50086 800 50194 856
rect 50362 800 50470 856
rect 50638 800 50746 856
rect 50914 800 51022 856
rect 51190 800 51298 856
rect 51466 800 51574 856
rect 51742 800 51850 856
rect 52018 800 52126 856
rect 52294 800 52402 856
rect 52570 800 52678 856
rect 52846 800 52954 856
rect 53122 800 53230 856
rect 53398 800 53506 856
rect 53674 800 53782 856
rect 53950 800 54058 856
rect 54226 800 54334 856
rect 54502 800 54610 856
rect 54778 800 54886 856
rect 55054 800 55162 856
rect 55330 800 55438 856
rect 55606 800 55714 856
rect 55882 800 55990 856
rect 56158 800 56266 856
rect 56434 800 56542 856
rect 56710 800 56818 856
rect 56986 800 57094 856
rect 57262 800 57370 856
rect 57538 800 57646 856
rect 57814 800 57922 856
rect 58090 800 58198 856
rect 58366 800 58474 856
rect 58642 800 58750 856
rect 58918 800 59026 856
rect 59194 800 59302 856
rect 59470 800 59578 856
rect 59746 800 59854 856
rect 60022 800 60130 856
rect 60298 800 60406 856
rect 60574 800 60682 856
rect 60850 800 60958 856
rect 61126 800 61234 856
rect 61402 800 61510 856
rect 61678 800 61786 856
rect 61954 800 62062 856
rect 62230 800 62338 856
rect 62506 800 62614 856
rect 62782 800 62890 856
rect 63058 800 63166 856
rect 63334 800 63442 856
rect 63610 800 63718 856
rect 63886 800 63994 856
rect 64162 800 64270 856
rect 64438 800 64546 856
rect 64714 800 64822 856
rect 64990 800 65098 856
rect 65266 800 65374 856
rect 65542 800 65650 856
rect 65818 800 65926 856
rect 66094 800 66202 856
rect 66370 800 66478 856
rect 66646 800 66754 856
rect 66922 800 67030 856
rect 67198 800 67306 856
rect 67474 800 67582 856
rect 67750 800 67858 856
rect 68026 800 68134 856
rect 68302 800 68410 856
rect 68578 800 68686 856
rect 68854 800 68962 856
rect 69130 800 69238 856
rect 69406 800 69514 856
rect 69682 800 69790 856
rect 69958 800 70066 856
rect 70234 800 70342 856
rect 70510 800 70618 856
rect 70786 800 70894 856
rect 71062 800 71170 856
rect 71338 800 71446 856
rect 71614 800 71722 856
rect 71890 800 71998 856
rect 72166 800 72274 856
rect 72442 800 72550 856
rect 72718 800 72826 856
rect 72994 800 73102 856
rect 73270 800 73378 856
rect 73546 800 73654 856
rect 73822 800 73930 856
rect 74098 800 74206 856
rect 74374 800 74482 856
rect 74650 800 74758 856
rect 74926 800 75034 856
rect 75202 800 75310 856
rect 75478 800 75586 856
rect 75754 800 75862 856
rect 76030 800 76138 856
rect 76306 800 76414 856
rect 76582 800 76690 856
rect 76858 800 76966 856
rect 77134 800 77242 856
rect 77410 800 77518 856
rect 77686 800 77794 856
rect 77962 800 78070 856
rect 78238 800 78346 856
rect 78514 800 78622 856
rect 78790 800 78898 856
rect 79066 800 79174 856
rect 79342 800 79450 856
rect 79618 800 79726 856
rect 79894 800 80002 856
rect 80170 800 80278 856
rect 80446 800 80554 856
rect 80722 800 80830 856
rect 80998 800 81106 856
rect 81274 800 81382 856
rect 81550 800 81658 856
rect 81826 800 81934 856
rect 82102 800 82210 856
rect 82378 800 82486 856
rect 82654 800 82762 856
rect 82930 800 83038 856
rect 83206 800 83314 856
rect 83482 800 83590 856
rect 83758 800 83866 856
rect 84034 800 84142 856
rect 84310 800 84418 856
rect 84586 800 84694 856
rect 84862 800 84970 856
rect 85138 800 85246 856
rect 85414 800 85522 856
rect 85690 800 85798 856
rect 85966 800 86074 856
rect 86242 800 86350 856
rect 86518 800 86626 856
rect 86794 800 86902 856
rect 87070 800 87178 856
rect 87346 800 87454 856
rect 87622 800 87730 856
rect 87898 800 88006 856
rect 88174 800 88282 856
rect 88450 800 88558 856
rect 88726 800 88834 856
rect 89002 800 89110 856
rect 89278 800 89386 856
rect 89554 800 89662 856
rect 89830 800 89938 856
rect 90106 800 90214 856
rect 90382 800 90490 856
rect 90658 800 90766 856
rect 90934 800 91042 856
rect 91210 800 91318 856
rect 91486 800 91594 856
rect 91762 800 91870 856
rect 92038 800 92146 856
rect 92314 800 92422 856
rect 92590 800 92698 856
rect 92866 800 92974 856
rect 93142 800 93250 856
rect 93418 800 93526 856
rect 93694 800 93802 856
rect 93970 800 94078 856
rect 94246 800 94354 856
rect 94522 800 94630 856
rect 94798 800 94906 856
rect 95074 800 95182 856
rect 95350 800 95458 856
rect 95626 800 95734 856
rect 95902 800 96010 856
rect 96178 800 96286 856
rect 96454 800 96562 856
rect 96730 800 96838 856
rect 97006 800 97114 856
rect 97282 800 97390 856
rect 97558 800 97666 856
rect 97834 800 97942 856
rect 98110 800 98218 856
rect 98386 800 98494 856
rect 98662 800 98770 856
rect 98938 800 99046 856
rect 99214 800 99322 856
rect 99490 800 99598 856
rect 99766 800 99874 856
rect 100042 800 100150 856
rect 100318 800 100426 856
rect 100594 800 100702 856
rect 100870 800 100978 856
rect 101146 800 101254 856
rect 101422 800 101530 856
rect 101698 800 101806 856
rect 101974 800 102082 856
rect 102250 800 102358 856
rect 102526 800 102634 856
rect 102802 800 102910 856
rect 103078 800 103186 856
rect 103354 800 103462 856
rect 103630 800 103738 856
rect 103906 800 104014 856
rect 104182 800 104290 856
rect 104458 800 104566 856
rect 104734 800 104842 856
rect 105010 800 105118 856
rect 105286 800 105394 856
rect 105562 800 105670 856
rect 105838 800 105946 856
rect 106114 800 106222 856
rect 106390 800 106498 856
rect 106666 800 106774 856
rect 106942 800 107050 856
rect 107218 800 107326 856
rect 107494 800 107602 856
rect 107770 800 107878 856
rect 108046 800 108154 856
rect 108322 800 108430 856
rect 108598 800 108706 856
rect 108874 800 108982 856
rect 109150 800 109258 856
rect 109426 800 109534 856
rect 109702 800 109810 856
rect 109978 800 110086 856
rect 110254 800 110362 856
rect 110530 800 110638 856
rect 110806 800 110914 856
rect 111082 800 111190 856
rect 111358 800 111466 856
rect 111634 800 111742 856
rect 111910 800 112018 856
rect 112186 800 112294 856
rect 112462 800 112570 856
rect 112738 800 112846 856
rect 113014 800 113122 856
rect 113290 800 113398 856
rect 113566 800 113674 856
rect 113842 800 113950 856
rect 114118 800 114226 856
rect 114394 800 114502 856
rect 114670 800 114778 856
rect 114946 800 115054 856
rect 115222 800 115330 856
rect 115498 800 115606 856
rect 115774 800 115882 856
rect 116050 800 116158 856
rect 116326 800 116434 856
rect 116602 800 116710 856
rect 116878 800 116986 856
rect 117154 800 117262 856
rect 117430 800 117538 856
rect 117706 800 117814 856
rect 117982 800 118090 856
rect 118258 800 118366 856
rect 118534 800 118642 856
rect 118810 800 118918 856
rect 119086 800 119194 856
rect 119362 800 119470 856
rect 119638 800 119746 856
rect 119914 800 120022 856
rect 120190 800 120298 856
rect 120466 800 120574 856
rect 120742 800 120850 856
rect 121018 800 121126 856
rect 121294 800 121402 856
rect 121570 800 121678 856
rect 121846 800 121954 856
rect 122122 800 122230 856
rect 122398 800 122506 856
rect 122674 800 122782 856
rect 122950 800 123058 856
rect 123226 800 123334 856
rect 123502 800 123610 856
rect 123778 800 123886 856
rect 124054 800 124162 856
rect 124330 800 124438 856
rect 124606 800 124714 856
rect 124882 800 124990 856
rect 125158 800 125266 856
rect 125434 800 125542 856
rect 125710 800 125818 856
rect 125986 800 126094 856
rect 126262 800 126370 856
rect 126538 800 126646 856
rect 126814 800 126922 856
rect 127090 800 127198 856
rect 127366 800 127474 856
rect 127642 800 127750 856
rect 127918 800 128026 856
rect 128194 800 128302 856
rect 128470 800 128578 856
rect 128746 800 128854 856
rect 129022 800 129130 856
rect 129298 800 129406 856
rect 129574 800 129682 856
rect 129850 800 129958 856
rect 130126 800 130234 856
rect 130402 800 130510 856
rect 130678 800 130786 856
rect 130954 800 131062 856
rect 131230 800 131338 856
rect 131506 800 131614 856
rect 131782 800 131890 856
rect 132058 800 132166 856
rect 132334 800 132442 856
rect 132610 800 132718 856
rect 132886 800 132994 856
rect 133162 800 133270 856
rect 133438 800 133546 856
rect 133714 800 133822 856
rect 133990 800 134098 856
rect 134266 800 134374 856
rect 134542 800 134650 856
rect 134818 800 134926 856
rect 135094 800 135202 856
rect 135370 800 135478 856
rect 135646 800 135754 856
rect 135922 800 136030 856
rect 136198 800 136306 856
rect 136474 800 136582 856
rect 136750 800 136858 856
rect 137026 800 137134 856
rect 137302 800 137410 856
rect 137578 800 137686 856
rect 137854 800 137962 856
rect 138130 800 138238 856
rect 138406 800 138514 856
rect 138682 800 138790 856
rect 138958 800 139066 856
rect 139234 800 139342 856
rect 139510 800 139618 856
rect 139786 800 139894 856
rect 140062 800 140170 856
rect 140338 800 140446 856
rect 140614 800 140722 856
rect 140890 800 140998 856
rect 141166 800 141274 856
rect 141442 800 141550 856
rect 141718 800 141826 856
rect 141994 800 142102 856
rect 142270 800 142378 856
rect 142546 800 142654 856
rect 142822 800 142930 856
rect 143098 800 143206 856
rect 143374 800 143482 856
rect 143650 800 143758 856
rect 143926 800 144034 856
rect 144202 800 144310 856
rect 144478 800 144586 856
rect 144754 800 144862 856
rect 145030 800 145138 856
rect 145306 800 145414 856
rect 145582 800 145690 856
rect 145858 800 145966 856
rect 146134 800 146242 856
rect 146410 800 146518 856
rect 146686 800 146794 856
rect 146962 800 147070 856
rect 147238 800 147346 856
rect 147514 800 147622 856
rect 147790 800 147898 856
rect 148066 800 159050 856
<< metal3 >>
rect 159200 157632 160000 157752
rect 0 155592 800 155712
rect 159200 154640 160000 154760
rect 0 152736 800 152856
rect 159200 151648 160000 151768
rect 0 149880 800 150000
rect 159200 148656 160000 148776
rect 0 147024 800 147144
rect 159200 145664 160000 145784
rect 0 144168 800 144288
rect 159200 142672 160000 142792
rect 0 141312 800 141432
rect 159200 139680 160000 139800
rect 0 138456 800 138576
rect 159200 136688 160000 136808
rect 0 135600 800 135720
rect 159200 133696 160000 133816
rect 0 132744 800 132864
rect 159200 130704 160000 130824
rect 0 129888 800 130008
rect 159200 127712 160000 127832
rect 0 127032 800 127152
rect 159200 124720 160000 124840
rect 0 124176 800 124296
rect 159200 121728 160000 121848
rect 0 121320 800 121440
rect 159200 118736 160000 118856
rect 0 118464 800 118584
rect 0 115608 800 115728
rect 159200 115744 160000 115864
rect 0 112752 800 112872
rect 159200 112752 160000 112872
rect 0 109896 800 110016
rect 159200 109760 160000 109880
rect 0 107040 800 107160
rect 159200 106768 160000 106888
rect 0 104184 800 104304
rect 159200 103776 160000 103896
rect 0 101328 800 101448
rect 159200 100784 160000 100904
rect 0 98472 800 98592
rect 159200 97792 160000 97912
rect 0 95616 800 95736
rect 159200 94800 160000 94920
rect 0 92760 800 92880
rect 159200 91808 160000 91928
rect 0 89904 800 90024
rect 159200 88816 160000 88936
rect 0 87048 800 87168
rect 159200 85824 160000 85944
rect 0 84192 800 84312
rect 159200 82832 160000 82952
rect 0 81336 800 81456
rect 159200 79840 160000 79960
rect 0 78480 800 78600
rect 159200 76848 160000 76968
rect 0 75624 800 75744
rect 159200 73856 160000 73976
rect 0 72768 800 72888
rect 159200 70864 160000 70984
rect 0 69912 800 70032
rect 159200 67872 160000 67992
rect 0 67056 800 67176
rect 159200 64880 160000 65000
rect 0 64200 800 64320
rect 159200 61888 160000 62008
rect 0 61344 800 61464
rect 159200 58896 160000 59016
rect 0 58488 800 58608
rect 159200 55904 160000 56024
rect 0 55632 800 55752
rect 0 52776 800 52896
rect 159200 52912 160000 53032
rect 0 49920 800 50040
rect 159200 49920 160000 50040
rect 0 47064 800 47184
rect 159200 46928 160000 47048
rect 0 44208 800 44328
rect 159200 43936 160000 44056
rect 0 41352 800 41472
rect 159200 40944 160000 41064
rect 0 38496 800 38616
rect 159200 37952 160000 38072
rect 0 35640 800 35760
rect 159200 34960 160000 35080
rect 0 32784 800 32904
rect 159200 31968 160000 32088
rect 0 29928 800 30048
rect 159200 28976 160000 29096
rect 0 27072 800 27192
rect 159200 25984 160000 26104
rect 0 24216 800 24336
rect 159200 22992 160000 23112
rect 0 21360 800 21480
rect 159200 20000 160000 20120
rect 0 18504 800 18624
rect 159200 17008 160000 17128
rect 0 15648 800 15768
rect 159200 14016 160000 14136
rect 0 12792 800 12912
rect 159200 11024 160000 11144
rect 0 9936 800 10056
rect 159200 8032 160000 8152
rect 0 7080 800 7200
rect 159200 5040 160000 5160
rect 0 4224 800 4344
rect 159200 2048 160000 2168
<< obsm3 >>
rect 800 157552 159120 157793
rect 800 155792 159200 157552
rect 880 155512 159200 155792
rect 800 154840 159200 155512
rect 800 154560 159120 154840
rect 800 152936 159200 154560
rect 880 152656 159200 152936
rect 800 151848 159200 152656
rect 800 151568 159120 151848
rect 800 150080 159200 151568
rect 880 149800 159200 150080
rect 800 148856 159200 149800
rect 800 148576 159120 148856
rect 800 147224 159200 148576
rect 880 146944 159200 147224
rect 800 145864 159200 146944
rect 800 145584 159120 145864
rect 800 144368 159200 145584
rect 880 144088 159200 144368
rect 800 142872 159200 144088
rect 800 142592 159120 142872
rect 800 141512 159200 142592
rect 880 141232 159200 141512
rect 800 139880 159200 141232
rect 800 139600 159120 139880
rect 800 138656 159200 139600
rect 880 138376 159200 138656
rect 800 136888 159200 138376
rect 800 136608 159120 136888
rect 800 135800 159200 136608
rect 880 135520 159200 135800
rect 800 133896 159200 135520
rect 800 133616 159120 133896
rect 800 132944 159200 133616
rect 880 132664 159200 132944
rect 800 130904 159200 132664
rect 800 130624 159120 130904
rect 800 130088 159200 130624
rect 880 129808 159200 130088
rect 800 127912 159200 129808
rect 800 127632 159120 127912
rect 800 127232 159200 127632
rect 880 126952 159200 127232
rect 800 124920 159200 126952
rect 800 124640 159120 124920
rect 800 124376 159200 124640
rect 880 124096 159200 124376
rect 800 121928 159200 124096
rect 800 121648 159120 121928
rect 800 121520 159200 121648
rect 880 121240 159200 121520
rect 800 118936 159200 121240
rect 800 118664 159120 118936
rect 880 118656 159120 118664
rect 880 118384 159200 118656
rect 800 115944 159200 118384
rect 800 115808 159120 115944
rect 880 115664 159120 115808
rect 880 115528 159200 115664
rect 800 112952 159200 115528
rect 880 112672 159120 112952
rect 800 110096 159200 112672
rect 880 109960 159200 110096
rect 880 109816 159120 109960
rect 800 109680 159120 109816
rect 800 107240 159200 109680
rect 880 106968 159200 107240
rect 880 106960 159120 106968
rect 800 106688 159120 106960
rect 800 104384 159200 106688
rect 880 104104 159200 104384
rect 800 103976 159200 104104
rect 800 103696 159120 103976
rect 800 101528 159200 103696
rect 880 101248 159200 101528
rect 800 100984 159200 101248
rect 800 100704 159120 100984
rect 800 98672 159200 100704
rect 880 98392 159200 98672
rect 800 97992 159200 98392
rect 800 97712 159120 97992
rect 800 95816 159200 97712
rect 880 95536 159200 95816
rect 800 95000 159200 95536
rect 800 94720 159120 95000
rect 800 92960 159200 94720
rect 880 92680 159200 92960
rect 800 92008 159200 92680
rect 800 91728 159120 92008
rect 800 90104 159200 91728
rect 880 89824 159200 90104
rect 800 89016 159200 89824
rect 800 88736 159120 89016
rect 800 87248 159200 88736
rect 880 86968 159200 87248
rect 800 86024 159200 86968
rect 800 85744 159120 86024
rect 800 84392 159200 85744
rect 880 84112 159200 84392
rect 800 83032 159200 84112
rect 800 82752 159120 83032
rect 800 81536 159200 82752
rect 880 81256 159200 81536
rect 800 80040 159200 81256
rect 800 79760 159120 80040
rect 800 78680 159200 79760
rect 880 78400 159200 78680
rect 800 77048 159200 78400
rect 800 76768 159120 77048
rect 800 75824 159200 76768
rect 880 75544 159200 75824
rect 800 74056 159200 75544
rect 800 73776 159120 74056
rect 800 72968 159200 73776
rect 880 72688 159200 72968
rect 800 71064 159200 72688
rect 800 70784 159120 71064
rect 800 70112 159200 70784
rect 880 69832 159200 70112
rect 800 68072 159200 69832
rect 800 67792 159120 68072
rect 800 67256 159200 67792
rect 880 66976 159200 67256
rect 800 65080 159200 66976
rect 800 64800 159120 65080
rect 800 64400 159200 64800
rect 880 64120 159200 64400
rect 800 62088 159200 64120
rect 800 61808 159120 62088
rect 800 61544 159200 61808
rect 880 61264 159200 61544
rect 800 59096 159200 61264
rect 800 58816 159120 59096
rect 800 58688 159200 58816
rect 880 58408 159200 58688
rect 800 56104 159200 58408
rect 800 55832 159120 56104
rect 880 55824 159120 55832
rect 880 55552 159200 55824
rect 800 53112 159200 55552
rect 800 52976 159120 53112
rect 880 52832 159120 52976
rect 880 52696 159200 52832
rect 800 50120 159200 52696
rect 880 49840 159120 50120
rect 800 47264 159200 49840
rect 880 47128 159200 47264
rect 880 46984 159120 47128
rect 800 46848 159120 46984
rect 800 44408 159200 46848
rect 880 44136 159200 44408
rect 880 44128 159120 44136
rect 800 43856 159120 44128
rect 800 41552 159200 43856
rect 880 41272 159200 41552
rect 800 41144 159200 41272
rect 800 40864 159120 41144
rect 800 38696 159200 40864
rect 880 38416 159200 38696
rect 800 38152 159200 38416
rect 800 37872 159120 38152
rect 800 35840 159200 37872
rect 880 35560 159200 35840
rect 800 35160 159200 35560
rect 800 34880 159120 35160
rect 800 32984 159200 34880
rect 880 32704 159200 32984
rect 800 32168 159200 32704
rect 800 31888 159120 32168
rect 800 30128 159200 31888
rect 880 29848 159200 30128
rect 800 29176 159200 29848
rect 800 28896 159120 29176
rect 800 27272 159200 28896
rect 880 26992 159200 27272
rect 800 26184 159200 26992
rect 800 25904 159120 26184
rect 800 24416 159200 25904
rect 880 24136 159200 24416
rect 800 23192 159200 24136
rect 800 22912 159120 23192
rect 800 21560 159200 22912
rect 880 21280 159200 21560
rect 800 20200 159200 21280
rect 800 19920 159120 20200
rect 800 18704 159200 19920
rect 880 18424 159200 18704
rect 800 17208 159200 18424
rect 800 16928 159120 17208
rect 800 15848 159200 16928
rect 880 15568 159200 15848
rect 800 14216 159200 15568
rect 800 13936 159120 14216
rect 800 12992 159200 13936
rect 880 12712 159200 12992
rect 800 11224 159200 12712
rect 800 10944 159120 11224
rect 800 10136 159200 10944
rect 880 9856 159200 10136
rect 800 8232 159200 9856
rect 800 7952 159120 8232
rect 800 7280 159200 7952
rect 880 7000 159200 7280
rect 800 5240 159200 7000
rect 800 4960 159120 5240
rect 800 4424 159200 4960
rect 880 4144 159200 4424
rect 800 2248 159200 4144
rect 800 2075 159120 2248
<< metal4 >>
rect 4208 2128 4528 157808
rect 4868 2128 5188 157808
rect 34928 2128 35248 157808
rect 35588 2128 35908 157808
rect 65648 2128 65968 157808
rect 66308 2128 66628 157808
rect 96368 2128 96688 157808
rect 97028 2128 97348 157808
rect 127088 2128 127408 157808
rect 127748 2128 128068 157808
rect 157808 2128 158128 157808
rect 158468 2128 158788 157808
<< obsm4 >>
rect 124811 56475 127008 149837
rect 127488 56475 127668 149837
rect 128148 56475 157261 149837
<< metal5 >>
rect 1056 128550 158932 128870
rect 1056 127890 158932 128210
rect 1056 97914 158932 98234
rect 1056 97254 158932 97574
rect 1056 67278 158932 67598
rect 1056 66618 158932 66938
rect 1056 36642 158932 36962
rect 1056 35982 158932 36302
rect 1056 6006 158932 6326
rect 1056 5346 158932 5666
<< labels >>
rlabel metal4 s 4868 2128 5188 157808 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 35588 2128 35908 157808 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 66308 2128 66628 157808 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 97028 2128 97348 157808 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127748 2128 128068 157808 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 158468 2128 158788 157808 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 6006 158932 6326 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 36642 158932 36962 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 67278 158932 67598 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 97914 158932 98234 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 128550 158932 128870 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 157808 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 157808 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 157808 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 157808 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 157808 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 157808 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5346 158932 5666 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 35982 158932 36302 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 66618 158932 66938 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 97254 158932 97574 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 127890 158932 128210 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 159200 64880 160000 65000 6 analog_io[0]
port 3 nsew signal bidirectional
rlabel metal2 s 121918 159200 121974 160000 6 analog_io[10]
port 4 nsew signal bidirectional
rlabel metal2 s 104254 159200 104310 160000 6 analog_io[11]
port 5 nsew signal bidirectional
rlabel metal2 s 86590 159200 86646 160000 6 analog_io[12]
port 6 nsew signal bidirectional
rlabel metal2 s 68926 159200 68982 160000 6 analog_io[13]
port 7 nsew signal bidirectional
rlabel metal2 s 51262 159200 51318 160000 6 analog_io[14]
port 8 nsew signal bidirectional
rlabel metal2 s 33598 159200 33654 160000 6 analog_io[15]
port 9 nsew signal bidirectional
rlabel metal2 s 15934 159200 15990 160000 6 analog_io[16]
port 10 nsew signal bidirectional
rlabel metal3 s 0 155592 800 155712 6 analog_io[17]
port 11 nsew signal bidirectional
rlabel metal3 s 0 144168 800 144288 6 analog_io[18]
port 12 nsew signal bidirectional
rlabel metal3 s 0 132744 800 132864 6 analog_io[19]
port 13 nsew signal bidirectional
rlabel metal3 s 159200 76848 160000 76968 6 analog_io[1]
port 14 nsew signal bidirectional
rlabel metal3 s 0 121320 800 121440 6 analog_io[20]
port 15 nsew signal bidirectional
rlabel metal3 s 0 109896 800 110016 6 analog_io[21]
port 16 nsew signal bidirectional
rlabel metal3 s 0 98472 800 98592 6 analog_io[22]
port 17 nsew signal bidirectional
rlabel metal3 s 0 87048 800 87168 6 analog_io[23]
port 18 nsew signal bidirectional
rlabel metal3 s 0 75624 800 75744 6 analog_io[24]
port 19 nsew signal bidirectional
rlabel metal3 s 0 64200 800 64320 6 analog_io[25]
port 20 nsew signal bidirectional
rlabel metal3 s 0 52776 800 52896 6 analog_io[26]
port 21 nsew signal bidirectional
rlabel metal3 s 0 41352 800 41472 6 analog_io[27]
port 22 nsew signal bidirectional
rlabel metal3 s 0 29928 800 30048 6 analog_io[28]
port 23 nsew signal bidirectional
rlabel metal3 s 159200 88816 160000 88936 6 analog_io[2]
port 24 nsew signal bidirectional
rlabel metal3 s 159200 100784 160000 100904 6 analog_io[3]
port 25 nsew signal bidirectional
rlabel metal3 s 159200 112752 160000 112872 6 analog_io[4]
port 26 nsew signal bidirectional
rlabel metal3 s 159200 124720 160000 124840 6 analog_io[5]
port 27 nsew signal bidirectional
rlabel metal3 s 159200 136688 160000 136808 6 analog_io[6]
port 28 nsew signal bidirectional
rlabel metal3 s 159200 148656 160000 148776 6 analog_io[7]
port 29 nsew signal bidirectional
rlabel metal2 s 157246 159200 157302 160000 6 analog_io[8]
port 30 nsew signal bidirectional
rlabel metal2 s 139582 159200 139638 160000 6 analog_io[9]
port 31 nsew signal bidirectional
rlabel metal3 s 159200 2048 160000 2168 6 io_in[0]
port 32 nsew signal input
rlabel metal3 s 159200 103776 160000 103896 6 io_in[10]
port 33 nsew signal input
rlabel metal3 s 159200 115744 160000 115864 6 io_in[11]
port 34 nsew signal input
rlabel metal3 s 159200 127712 160000 127832 6 io_in[12]
port 35 nsew signal input
rlabel metal3 s 159200 139680 160000 139800 6 io_in[13]
port 36 nsew signal input
rlabel metal3 s 159200 151648 160000 151768 6 io_in[14]
port 37 nsew signal input
rlabel metal2 s 152830 159200 152886 160000 6 io_in[15]
port 38 nsew signal input
rlabel metal2 s 135166 159200 135222 160000 6 io_in[16]
port 39 nsew signal input
rlabel metal2 s 117502 159200 117558 160000 6 io_in[17]
port 40 nsew signal input
rlabel metal2 s 99838 159200 99894 160000 6 io_in[18]
port 41 nsew signal input
rlabel metal2 s 82174 159200 82230 160000 6 io_in[19]
port 42 nsew signal input
rlabel metal3 s 159200 11024 160000 11144 6 io_in[1]
port 43 nsew signal input
rlabel metal2 s 64510 159200 64566 160000 6 io_in[20]
port 44 nsew signal input
rlabel metal2 s 46846 159200 46902 160000 6 io_in[21]
port 45 nsew signal input
rlabel metal2 s 29182 159200 29238 160000 6 io_in[22]
port 46 nsew signal input
rlabel metal2 s 11518 159200 11574 160000 6 io_in[23]
port 47 nsew signal input
rlabel metal3 s 0 152736 800 152856 6 io_in[24]
port 48 nsew signal input
rlabel metal3 s 0 141312 800 141432 6 io_in[25]
port 49 nsew signal input
rlabel metal3 s 0 129888 800 130008 6 io_in[26]
port 50 nsew signal input
rlabel metal3 s 0 118464 800 118584 6 io_in[27]
port 51 nsew signal input
rlabel metal3 s 0 107040 800 107160 6 io_in[28]
port 52 nsew signal input
rlabel metal3 s 0 95616 800 95736 6 io_in[29]
port 53 nsew signal input
rlabel metal3 s 159200 20000 160000 20120 6 io_in[2]
port 54 nsew signal input
rlabel metal3 s 0 84192 800 84312 6 io_in[30]
port 55 nsew signal input
rlabel metal3 s 0 72768 800 72888 6 io_in[31]
port 56 nsew signal input
rlabel metal3 s 0 61344 800 61464 6 io_in[32]
port 57 nsew signal input
rlabel metal3 s 0 49920 800 50040 6 io_in[33]
port 58 nsew signal input
rlabel metal3 s 0 38496 800 38616 6 io_in[34]
port 59 nsew signal input
rlabel metal3 s 0 27072 800 27192 6 io_in[35]
port 60 nsew signal input
rlabel metal3 s 0 18504 800 18624 6 io_in[36]
port 61 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 io_in[37]
port 62 nsew signal input
rlabel metal3 s 159200 28976 160000 29096 6 io_in[3]
port 63 nsew signal input
rlabel metal3 s 159200 37952 160000 38072 6 io_in[4]
port 64 nsew signal input
rlabel metal3 s 159200 46928 160000 47048 6 io_in[5]
port 65 nsew signal input
rlabel metal3 s 159200 55904 160000 56024 6 io_in[6]
port 66 nsew signal input
rlabel metal3 s 159200 67872 160000 67992 6 io_in[7]
port 67 nsew signal input
rlabel metal3 s 159200 79840 160000 79960 6 io_in[8]
port 68 nsew signal input
rlabel metal3 s 159200 91808 160000 91928 6 io_in[9]
port 69 nsew signal input
rlabel metal3 s 159200 8032 160000 8152 6 io_oeb[0]
port 70 nsew signal output
rlabel metal3 s 159200 109760 160000 109880 6 io_oeb[10]
port 71 nsew signal output
rlabel metal3 s 159200 121728 160000 121848 6 io_oeb[11]
port 72 nsew signal output
rlabel metal3 s 159200 133696 160000 133816 6 io_oeb[12]
port 73 nsew signal output
rlabel metal3 s 159200 145664 160000 145784 6 io_oeb[13]
port 74 nsew signal output
rlabel metal3 s 159200 157632 160000 157752 6 io_oeb[14]
port 75 nsew signal output
rlabel metal2 s 143998 159200 144054 160000 6 io_oeb[15]
port 76 nsew signal output
rlabel metal2 s 126334 159200 126390 160000 6 io_oeb[16]
port 77 nsew signal output
rlabel metal2 s 108670 159200 108726 160000 6 io_oeb[17]
port 78 nsew signal output
rlabel metal2 s 91006 159200 91062 160000 6 io_oeb[18]
port 79 nsew signal output
rlabel metal2 s 73342 159200 73398 160000 6 io_oeb[19]
port 80 nsew signal output
rlabel metal3 s 159200 17008 160000 17128 6 io_oeb[1]
port 81 nsew signal output
rlabel metal2 s 55678 159200 55734 160000 6 io_oeb[20]
port 82 nsew signal output
rlabel metal2 s 38014 159200 38070 160000 6 io_oeb[21]
port 83 nsew signal output
rlabel metal2 s 20350 159200 20406 160000 6 io_oeb[22]
port 84 nsew signal output
rlabel metal2 s 2686 159200 2742 160000 6 io_oeb[23]
port 85 nsew signal output
rlabel metal3 s 0 147024 800 147144 6 io_oeb[24]
port 86 nsew signal output
rlabel metal3 s 0 135600 800 135720 6 io_oeb[25]
port 87 nsew signal output
rlabel metal3 s 0 124176 800 124296 6 io_oeb[26]
port 88 nsew signal output
rlabel metal3 s 0 112752 800 112872 6 io_oeb[27]
port 89 nsew signal output
rlabel metal3 s 0 101328 800 101448 6 io_oeb[28]
port 90 nsew signal output
rlabel metal3 s 0 89904 800 90024 6 io_oeb[29]
port 91 nsew signal output
rlabel metal3 s 159200 25984 160000 26104 6 io_oeb[2]
port 92 nsew signal output
rlabel metal3 s 0 78480 800 78600 6 io_oeb[30]
port 93 nsew signal output
rlabel metal3 s 0 67056 800 67176 6 io_oeb[31]
port 94 nsew signal output
rlabel metal3 s 0 55632 800 55752 6 io_oeb[32]
port 95 nsew signal output
rlabel metal3 s 0 44208 800 44328 6 io_oeb[33]
port 96 nsew signal output
rlabel metal3 s 0 32784 800 32904 6 io_oeb[34]
port 97 nsew signal output
rlabel metal3 s 0 21360 800 21480 6 io_oeb[35]
port 98 nsew signal output
rlabel metal3 s 0 12792 800 12912 6 io_oeb[36]
port 99 nsew signal output
rlabel metal3 s 0 4224 800 4344 6 io_oeb[37]
port 100 nsew signal output
rlabel metal3 s 159200 34960 160000 35080 6 io_oeb[3]
port 101 nsew signal output
rlabel metal3 s 159200 43936 160000 44056 6 io_oeb[4]
port 102 nsew signal output
rlabel metal3 s 159200 52912 160000 53032 6 io_oeb[5]
port 103 nsew signal output
rlabel metal3 s 159200 61888 160000 62008 6 io_oeb[6]
port 104 nsew signal output
rlabel metal3 s 159200 73856 160000 73976 6 io_oeb[7]
port 105 nsew signal output
rlabel metal3 s 159200 85824 160000 85944 6 io_oeb[8]
port 106 nsew signal output
rlabel metal3 s 159200 97792 160000 97912 6 io_oeb[9]
port 107 nsew signal output
rlabel metal3 s 159200 5040 160000 5160 6 io_out[0]
port 108 nsew signal output
rlabel metal3 s 159200 106768 160000 106888 6 io_out[10]
port 109 nsew signal output
rlabel metal3 s 159200 118736 160000 118856 6 io_out[11]
port 110 nsew signal output
rlabel metal3 s 159200 130704 160000 130824 6 io_out[12]
port 111 nsew signal output
rlabel metal3 s 159200 142672 160000 142792 6 io_out[13]
port 112 nsew signal output
rlabel metal3 s 159200 154640 160000 154760 6 io_out[14]
port 113 nsew signal output
rlabel metal2 s 148414 159200 148470 160000 6 io_out[15]
port 114 nsew signal output
rlabel metal2 s 130750 159200 130806 160000 6 io_out[16]
port 115 nsew signal output
rlabel metal2 s 113086 159200 113142 160000 6 io_out[17]
port 116 nsew signal output
rlabel metal2 s 95422 159200 95478 160000 6 io_out[18]
port 117 nsew signal output
rlabel metal2 s 77758 159200 77814 160000 6 io_out[19]
port 118 nsew signal output
rlabel metal3 s 159200 14016 160000 14136 6 io_out[1]
port 119 nsew signal output
rlabel metal2 s 60094 159200 60150 160000 6 io_out[20]
port 120 nsew signal output
rlabel metal2 s 42430 159200 42486 160000 6 io_out[21]
port 121 nsew signal output
rlabel metal2 s 24766 159200 24822 160000 6 io_out[22]
port 122 nsew signal output
rlabel metal2 s 7102 159200 7158 160000 6 io_out[23]
port 123 nsew signal output
rlabel metal3 s 0 149880 800 150000 6 io_out[24]
port 124 nsew signal output
rlabel metal3 s 0 138456 800 138576 6 io_out[25]
port 125 nsew signal output
rlabel metal3 s 0 127032 800 127152 6 io_out[26]
port 126 nsew signal output
rlabel metal3 s 0 115608 800 115728 6 io_out[27]
port 127 nsew signal output
rlabel metal3 s 0 104184 800 104304 6 io_out[28]
port 128 nsew signal output
rlabel metal3 s 0 92760 800 92880 6 io_out[29]
port 129 nsew signal output
rlabel metal3 s 159200 22992 160000 23112 6 io_out[2]
port 130 nsew signal output
rlabel metal3 s 0 81336 800 81456 6 io_out[30]
port 131 nsew signal output
rlabel metal3 s 0 69912 800 70032 6 io_out[31]
port 132 nsew signal output
rlabel metal3 s 0 58488 800 58608 6 io_out[32]
port 133 nsew signal output
rlabel metal3 s 0 47064 800 47184 6 io_out[33]
port 134 nsew signal output
rlabel metal3 s 0 35640 800 35760 6 io_out[34]
port 135 nsew signal output
rlabel metal3 s 0 24216 800 24336 6 io_out[35]
port 136 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 io_out[36]
port 137 nsew signal output
rlabel metal3 s 0 7080 800 7200 6 io_out[37]
port 138 nsew signal output
rlabel metal3 s 159200 31968 160000 32088 6 io_out[3]
port 139 nsew signal output
rlabel metal3 s 159200 40944 160000 41064 6 io_out[4]
port 140 nsew signal output
rlabel metal3 s 159200 49920 160000 50040 6 io_out[5]
port 141 nsew signal output
rlabel metal3 s 159200 58896 160000 59016 6 io_out[6]
port 142 nsew signal output
rlabel metal3 s 159200 70864 160000 70984 6 io_out[7]
port 143 nsew signal output
rlabel metal3 s 159200 82832 160000 82952 6 io_out[8]
port 144 nsew signal output
rlabel metal3 s 159200 94800 160000 94920 6 io_out[9]
port 145 nsew signal output
rlabel metal2 s 41142 0 41198 800 6 la_data_in[0]
port 146 nsew signal input
rlabel metal2 s 123942 0 123998 800 6 la_data_in[100]
port 147 nsew signal input
rlabel metal2 s 124770 0 124826 800 6 la_data_in[101]
port 148 nsew signal input
rlabel metal2 s 125598 0 125654 800 6 la_data_in[102]
port 149 nsew signal input
rlabel metal2 s 126426 0 126482 800 6 la_data_in[103]
port 150 nsew signal input
rlabel metal2 s 127254 0 127310 800 6 la_data_in[104]
port 151 nsew signal input
rlabel metal2 s 128082 0 128138 800 6 la_data_in[105]
port 152 nsew signal input
rlabel metal2 s 128910 0 128966 800 6 la_data_in[106]
port 153 nsew signal input
rlabel metal2 s 129738 0 129794 800 6 la_data_in[107]
port 154 nsew signal input
rlabel metal2 s 130566 0 130622 800 6 la_data_in[108]
port 155 nsew signal input
rlabel metal2 s 131394 0 131450 800 6 la_data_in[109]
port 156 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 la_data_in[10]
port 157 nsew signal input
rlabel metal2 s 132222 0 132278 800 6 la_data_in[110]
port 158 nsew signal input
rlabel metal2 s 133050 0 133106 800 6 la_data_in[111]
port 159 nsew signal input
rlabel metal2 s 133878 0 133934 800 6 la_data_in[112]
port 160 nsew signal input
rlabel metal2 s 134706 0 134762 800 6 la_data_in[113]
port 161 nsew signal input
rlabel metal2 s 135534 0 135590 800 6 la_data_in[114]
port 162 nsew signal input
rlabel metal2 s 136362 0 136418 800 6 la_data_in[115]
port 163 nsew signal input
rlabel metal2 s 137190 0 137246 800 6 la_data_in[116]
port 164 nsew signal input
rlabel metal2 s 138018 0 138074 800 6 la_data_in[117]
port 165 nsew signal input
rlabel metal2 s 138846 0 138902 800 6 la_data_in[118]
port 166 nsew signal input
rlabel metal2 s 139674 0 139730 800 6 la_data_in[119]
port 167 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 la_data_in[11]
port 168 nsew signal input
rlabel metal2 s 140502 0 140558 800 6 la_data_in[120]
port 169 nsew signal input
rlabel metal2 s 141330 0 141386 800 6 la_data_in[121]
port 170 nsew signal input
rlabel metal2 s 142158 0 142214 800 6 la_data_in[122]
port 171 nsew signal input
rlabel metal2 s 142986 0 143042 800 6 la_data_in[123]
port 172 nsew signal input
rlabel metal2 s 143814 0 143870 800 6 la_data_in[124]
port 173 nsew signal input
rlabel metal2 s 144642 0 144698 800 6 la_data_in[125]
port 174 nsew signal input
rlabel metal2 s 145470 0 145526 800 6 la_data_in[126]
port 175 nsew signal input
rlabel metal2 s 146298 0 146354 800 6 la_data_in[127]
port 176 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 la_data_in[12]
port 177 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 la_data_in[13]
port 178 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 la_data_in[14]
port 179 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 la_data_in[15]
port 180 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 la_data_in[16]
port 181 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 la_data_in[17]
port 182 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 la_data_in[18]
port 183 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 la_data_in[19]
port 184 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 la_data_in[1]
port 185 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 la_data_in[20]
port 186 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 la_data_in[21]
port 187 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 la_data_in[22]
port 188 nsew signal input
rlabel metal2 s 60186 0 60242 800 6 la_data_in[23]
port 189 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 la_data_in[24]
port 190 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 la_data_in[25]
port 191 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 la_data_in[26]
port 192 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 la_data_in[27]
port 193 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 la_data_in[28]
port 194 nsew signal input
rlabel metal2 s 65154 0 65210 800 6 la_data_in[29]
port 195 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 la_data_in[2]
port 196 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 la_data_in[30]
port 197 nsew signal input
rlabel metal2 s 66810 0 66866 800 6 la_data_in[31]
port 198 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 la_data_in[32]
port 199 nsew signal input
rlabel metal2 s 68466 0 68522 800 6 la_data_in[33]
port 200 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 la_data_in[34]
port 201 nsew signal input
rlabel metal2 s 70122 0 70178 800 6 la_data_in[35]
port 202 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 la_data_in[36]
port 203 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 la_data_in[37]
port 204 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 la_data_in[38]
port 205 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 la_data_in[39]
port 206 nsew signal input
rlabel metal2 s 43626 0 43682 800 6 la_data_in[3]
port 207 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 la_data_in[40]
port 208 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 la_data_in[41]
port 209 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 la_data_in[42]
port 210 nsew signal input
rlabel metal2 s 76746 0 76802 800 6 la_data_in[43]
port 211 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 la_data_in[44]
port 212 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 la_data_in[45]
port 213 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 la_data_in[46]
port 214 nsew signal input
rlabel metal2 s 80058 0 80114 800 6 la_data_in[47]
port 215 nsew signal input
rlabel metal2 s 80886 0 80942 800 6 la_data_in[48]
port 216 nsew signal input
rlabel metal2 s 81714 0 81770 800 6 la_data_in[49]
port 217 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 la_data_in[4]
port 218 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 la_data_in[50]
port 219 nsew signal input
rlabel metal2 s 83370 0 83426 800 6 la_data_in[51]
port 220 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 la_data_in[52]
port 221 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 la_data_in[53]
port 222 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 la_data_in[54]
port 223 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 la_data_in[55]
port 224 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 la_data_in[56]
port 225 nsew signal input
rlabel metal2 s 88338 0 88394 800 6 la_data_in[57]
port 226 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 la_data_in[58]
port 227 nsew signal input
rlabel metal2 s 89994 0 90050 800 6 la_data_in[59]
port 228 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 la_data_in[5]
port 229 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 la_data_in[60]
port 230 nsew signal input
rlabel metal2 s 91650 0 91706 800 6 la_data_in[61]
port 231 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 la_data_in[62]
port 232 nsew signal input
rlabel metal2 s 93306 0 93362 800 6 la_data_in[63]
port 233 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 la_data_in[64]
port 234 nsew signal input
rlabel metal2 s 94962 0 95018 800 6 la_data_in[65]
port 235 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_data_in[66]
port 236 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 la_data_in[67]
port 237 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_data_in[68]
port 238 nsew signal input
rlabel metal2 s 98274 0 98330 800 6 la_data_in[69]
port 239 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 la_data_in[6]
port 240 nsew signal input
rlabel metal2 s 99102 0 99158 800 6 la_data_in[70]
port 241 nsew signal input
rlabel metal2 s 99930 0 99986 800 6 la_data_in[71]
port 242 nsew signal input
rlabel metal2 s 100758 0 100814 800 6 la_data_in[72]
port 243 nsew signal input
rlabel metal2 s 101586 0 101642 800 6 la_data_in[73]
port 244 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 la_data_in[74]
port 245 nsew signal input
rlabel metal2 s 103242 0 103298 800 6 la_data_in[75]
port 246 nsew signal input
rlabel metal2 s 104070 0 104126 800 6 la_data_in[76]
port 247 nsew signal input
rlabel metal2 s 104898 0 104954 800 6 la_data_in[77]
port 248 nsew signal input
rlabel metal2 s 105726 0 105782 800 6 la_data_in[78]
port 249 nsew signal input
rlabel metal2 s 106554 0 106610 800 6 la_data_in[79]
port 250 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 la_data_in[7]
port 251 nsew signal input
rlabel metal2 s 107382 0 107438 800 6 la_data_in[80]
port 252 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 la_data_in[81]
port 253 nsew signal input
rlabel metal2 s 109038 0 109094 800 6 la_data_in[82]
port 254 nsew signal input
rlabel metal2 s 109866 0 109922 800 6 la_data_in[83]
port 255 nsew signal input
rlabel metal2 s 110694 0 110750 800 6 la_data_in[84]
port 256 nsew signal input
rlabel metal2 s 111522 0 111578 800 6 la_data_in[85]
port 257 nsew signal input
rlabel metal2 s 112350 0 112406 800 6 la_data_in[86]
port 258 nsew signal input
rlabel metal2 s 113178 0 113234 800 6 la_data_in[87]
port 259 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 la_data_in[88]
port 260 nsew signal input
rlabel metal2 s 114834 0 114890 800 6 la_data_in[89]
port 261 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 la_data_in[8]
port 262 nsew signal input
rlabel metal2 s 115662 0 115718 800 6 la_data_in[90]
port 263 nsew signal input
rlabel metal2 s 116490 0 116546 800 6 la_data_in[91]
port 264 nsew signal input
rlabel metal2 s 117318 0 117374 800 6 la_data_in[92]
port 265 nsew signal input
rlabel metal2 s 118146 0 118202 800 6 la_data_in[93]
port 266 nsew signal input
rlabel metal2 s 118974 0 119030 800 6 la_data_in[94]
port 267 nsew signal input
rlabel metal2 s 119802 0 119858 800 6 la_data_in[95]
port 268 nsew signal input
rlabel metal2 s 120630 0 120686 800 6 la_data_in[96]
port 269 nsew signal input
rlabel metal2 s 121458 0 121514 800 6 la_data_in[97]
port 270 nsew signal input
rlabel metal2 s 122286 0 122342 800 6 la_data_in[98]
port 271 nsew signal input
rlabel metal2 s 123114 0 123170 800 6 la_data_in[99]
port 272 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 la_data_in[9]
port 273 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 la_data_out[0]
port 274 nsew signal output
rlabel metal2 s 124218 0 124274 800 6 la_data_out[100]
port 275 nsew signal output
rlabel metal2 s 125046 0 125102 800 6 la_data_out[101]
port 276 nsew signal output
rlabel metal2 s 125874 0 125930 800 6 la_data_out[102]
port 277 nsew signal output
rlabel metal2 s 126702 0 126758 800 6 la_data_out[103]
port 278 nsew signal output
rlabel metal2 s 127530 0 127586 800 6 la_data_out[104]
port 279 nsew signal output
rlabel metal2 s 128358 0 128414 800 6 la_data_out[105]
port 280 nsew signal output
rlabel metal2 s 129186 0 129242 800 6 la_data_out[106]
port 281 nsew signal output
rlabel metal2 s 130014 0 130070 800 6 la_data_out[107]
port 282 nsew signal output
rlabel metal2 s 130842 0 130898 800 6 la_data_out[108]
port 283 nsew signal output
rlabel metal2 s 131670 0 131726 800 6 la_data_out[109]
port 284 nsew signal output
rlabel metal2 s 49698 0 49754 800 6 la_data_out[10]
port 285 nsew signal output
rlabel metal2 s 132498 0 132554 800 6 la_data_out[110]
port 286 nsew signal output
rlabel metal2 s 133326 0 133382 800 6 la_data_out[111]
port 287 nsew signal output
rlabel metal2 s 134154 0 134210 800 6 la_data_out[112]
port 288 nsew signal output
rlabel metal2 s 134982 0 135038 800 6 la_data_out[113]
port 289 nsew signal output
rlabel metal2 s 135810 0 135866 800 6 la_data_out[114]
port 290 nsew signal output
rlabel metal2 s 136638 0 136694 800 6 la_data_out[115]
port 291 nsew signal output
rlabel metal2 s 137466 0 137522 800 6 la_data_out[116]
port 292 nsew signal output
rlabel metal2 s 138294 0 138350 800 6 la_data_out[117]
port 293 nsew signal output
rlabel metal2 s 139122 0 139178 800 6 la_data_out[118]
port 294 nsew signal output
rlabel metal2 s 139950 0 140006 800 6 la_data_out[119]
port 295 nsew signal output
rlabel metal2 s 50526 0 50582 800 6 la_data_out[11]
port 296 nsew signal output
rlabel metal2 s 140778 0 140834 800 6 la_data_out[120]
port 297 nsew signal output
rlabel metal2 s 141606 0 141662 800 6 la_data_out[121]
port 298 nsew signal output
rlabel metal2 s 142434 0 142490 800 6 la_data_out[122]
port 299 nsew signal output
rlabel metal2 s 143262 0 143318 800 6 la_data_out[123]
port 300 nsew signal output
rlabel metal2 s 144090 0 144146 800 6 la_data_out[124]
port 301 nsew signal output
rlabel metal2 s 144918 0 144974 800 6 la_data_out[125]
port 302 nsew signal output
rlabel metal2 s 145746 0 145802 800 6 la_data_out[126]
port 303 nsew signal output
rlabel metal2 s 146574 0 146630 800 6 la_data_out[127]
port 304 nsew signal output
rlabel metal2 s 51354 0 51410 800 6 la_data_out[12]
port 305 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 la_data_out[13]
port 306 nsew signal output
rlabel metal2 s 53010 0 53066 800 6 la_data_out[14]
port 307 nsew signal output
rlabel metal2 s 53838 0 53894 800 6 la_data_out[15]
port 308 nsew signal output
rlabel metal2 s 54666 0 54722 800 6 la_data_out[16]
port 309 nsew signal output
rlabel metal2 s 55494 0 55550 800 6 la_data_out[17]
port 310 nsew signal output
rlabel metal2 s 56322 0 56378 800 6 la_data_out[18]
port 311 nsew signal output
rlabel metal2 s 57150 0 57206 800 6 la_data_out[19]
port 312 nsew signal output
rlabel metal2 s 42246 0 42302 800 6 la_data_out[1]
port 313 nsew signal output
rlabel metal2 s 57978 0 58034 800 6 la_data_out[20]
port 314 nsew signal output
rlabel metal2 s 58806 0 58862 800 6 la_data_out[21]
port 315 nsew signal output
rlabel metal2 s 59634 0 59690 800 6 la_data_out[22]
port 316 nsew signal output
rlabel metal2 s 60462 0 60518 800 6 la_data_out[23]
port 317 nsew signal output
rlabel metal2 s 61290 0 61346 800 6 la_data_out[24]
port 318 nsew signal output
rlabel metal2 s 62118 0 62174 800 6 la_data_out[25]
port 319 nsew signal output
rlabel metal2 s 62946 0 63002 800 6 la_data_out[26]
port 320 nsew signal output
rlabel metal2 s 63774 0 63830 800 6 la_data_out[27]
port 321 nsew signal output
rlabel metal2 s 64602 0 64658 800 6 la_data_out[28]
port 322 nsew signal output
rlabel metal2 s 65430 0 65486 800 6 la_data_out[29]
port 323 nsew signal output
rlabel metal2 s 43074 0 43130 800 6 la_data_out[2]
port 324 nsew signal output
rlabel metal2 s 66258 0 66314 800 6 la_data_out[30]
port 325 nsew signal output
rlabel metal2 s 67086 0 67142 800 6 la_data_out[31]
port 326 nsew signal output
rlabel metal2 s 67914 0 67970 800 6 la_data_out[32]
port 327 nsew signal output
rlabel metal2 s 68742 0 68798 800 6 la_data_out[33]
port 328 nsew signal output
rlabel metal2 s 69570 0 69626 800 6 la_data_out[34]
port 329 nsew signal output
rlabel metal2 s 70398 0 70454 800 6 la_data_out[35]
port 330 nsew signal output
rlabel metal2 s 71226 0 71282 800 6 la_data_out[36]
port 331 nsew signal output
rlabel metal2 s 72054 0 72110 800 6 la_data_out[37]
port 332 nsew signal output
rlabel metal2 s 72882 0 72938 800 6 la_data_out[38]
port 333 nsew signal output
rlabel metal2 s 73710 0 73766 800 6 la_data_out[39]
port 334 nsew signal output
rlabel metal2 s 43902 0 43958 800 6 la_data_out[3]
port 335 nsew signal output
rlabel metal2 s 74538 0 74594 800 6 la_data_out[40]
port 336 nsew signal output
rlabel metal2 s 75366 0 75422 800 6 la_data_out[41]
port 337 nsew signal output
rlabel metal2 s 76194 0 76250 800 6 la_data_out[42]
port 338 nsew signal output
rlabel metal2 s 77022 0 77078 800 6 la_data_out[43]
port 339 nsew signal output
rlabel metal2 s 77850 0 77906 800 6 la_data_out[44]
port 340 nsew signal output
rlabel metal2 s 78678 0 78734 800 6 la_data_out[45]
port 341 nsew signal output
rlabel metal2 s 79506 0 79562 800 6 la_data_out[46]
port 342 nsew signal output
rlabel metal2 s 80334 0 80390 800 6 la_data_out[47]
port 343 nsew signal output
rlabel metal2 s 81162 0 81218 800 6 la_data_out[48]
port 344 nsew signal output
rlabel metal2 s 81990 0 82046 800 6 la_data_out[49]
port 345 nsew signal output
rlabel metal2 s 44730 0 44786 800 6 la_data_out[4]
port 346 nsew signal output
rlabel metal2 s 82818 0 82874 800 6 la_data_out[50]
port 347 nsew signal output
rlabel metal2 s 83646 0 83702 800 6 la_data_out[51]
port 348 nsew signal output
rlabel metal2 s 84474 0 84530 800 6 la_data_out[52]
port 349 nsew signal output
rlabel metal2 s 85302 0 85358 800 6 la_data_out[53]
port 350 nsew signal output
rlabel metal2 s 86130 0 86186 800 6 la_data_out[54]
port 351 nsew signal output
rlabel metal2 s 86958 0 87014 800 6 la_data_out[55]
port 352 nsew signal output
rlabel metal2 s 87786 0 87842 800 6 la_data_out[56]
port 353 nsew signal output
rlabel metal2 s 88614 0 88670 800 6 la_data_out[57]
port 354 nsew signal output
rlabel metal2 s 89442 0 89498 800 6 la_data_out[58]
port 355 nsew signal output
rlabel metal2 s 90270 0 90326 800 6 la_data_out[59]
port 356 nsew signal output
rlabel metal2 s 45558 0 45614 800 6 la_data_out[5]
port 357 nsew signal output
rlabel metal2 s 91098 0 91154 800 6 la_data_out[60]
port 358 nsew signal output
rlabel metal2 s 91926 0 91982 800 6 la_data_out[61]
port 359 nsew signal output
rlabel metal2 s 92754 0 92810 800 6 la_data_out[62]
port 360 nsew signal output
rlabel metal2 s 93582 0 93638 800 6 la_data_out[63]
port 361 nsew signal output
rlabel metal2 s 94410 0 94466 800 6 la_data_out[64]
port 362 nsew signal output
rlabel metal2 s 95238 0 95294 800 6 la_data_out[65]
port 363 nsew signal output
rlabel metal2 s 96066 0 96122 800 6 la_data_out[66]
port 364 nsew signal output
rlabel metal2 s 96894 0 96950 800 6 la_data_out[67]
port 365 nsew signal output
rlabel metal2 s 97722 0 97778 800 6 la_data_out[68]
port 366 nsew signal output
rlabel metal2 s 98550 0 98606 800 6 la_data_out[69]
port 367 nsew signal output
rlabel metal2 s 46386 0 46442 800 6 la_data_out[6]
port 368 nsew signal output
rlabel metal2 s 99378 0 99434 800 6 la_data_out[70]
port 369 nsew signal output
rlabel metal2 s 100206 0 100262 800 6 la_data_out[71]
port 370 nsew signal output
rlabel metal2 s 101034 0 101090 800 6 la_data_out[72]
port 371 nsew signal output
rlabel metal2 s 101862 0 101918 800 6 la_data_out[73]
port 372 nsew signal output
rlabel metal2 s 102690 0 102746 800 6 la_data_out[74]
port 373 nsew signal output
rlabel metal2 s 103518 0 103574 800 6 la_data_out[75]
port 374 nsew signal output
rlabel metal2 s 104346 0 104402 800 6 la_data_out[76]
port 375 nsew signal output
rlabel metal2 s 105174 0 105230 800 6 la_data_out[77]
port 376 nsew signal output
rlabel metal2 s 106002 0 106058 800 6 la_data_out[78]
port 377 nsew signal output
rlabel metal2 s 106830 0 106886 800 6 la_data_out[79]
port 378 nsew signal output
rlabel metal2 s 47214 0 47270 800 6 la_data_out[7]
port 379 nsew signal output
rlabel metal2 s 107658 0 107714 800 6 la_data_out[80]
port 380 nsew signal output
rlabel metal2 s 108486 0 108542 800 6 la_data_out[81]
port 381 nsew signal output
rlabel metal2 s 109314 0 109370 800 6 la_data_out[82]
port 382 nsew signal output
rlabel metal2 s 110142 0 110198 800 6 la_data_out[83]
port 383 nsew signal output
rlabel metal2 s 110970 0 111026 800 6 la_data_out[84]
port 384 nsew signal output
rlabel metal2 s 111798 0 111854 800 6 la_data_out[85]
port 385 nsew signal output
rlabel metal2 s 112626 0 112682 800 6 la_data_out[86]
port 386 nsew signal output
rlabel metal2 s 113454 0 113510 800 6 la_data_out[87]
port 387 nsew signal output
rlabel metal2 s 114282 0 114338 800 6 la_data_out[88]
port 388 nsew signal output
rlabel metal2 s 115110 0 115166 800 6 la_data_out[89]
port 389 nsew signal output
rlabel metal2 s 48042 0 48098 800 6 la_data_out[8]
port 390 nsew signal output
rlabel metal2 s 115938 0 115994 800 6 la_data_out[90]
port 391 nsew signal output
rlabel metal2 s 116766 0 116822 800 6 la_data_out[91]
port 392 nsew signal output
rlabel metal2 s 117594 0 117650 800 6 la_data_out[92]
port 393 nsew signal output
rlabel metal2 s 118422 0 118478 800 6 la_data_out[93]
port 394 nsew signal output
rlabel metal2 s 119250 0 119306 800 6 la_data_out[94]
port 395 nsew signal output
rlabel metal2 s 120078 0 120134 800 6 la_data_out[95]
port 396 nsew signal output
rlabel metal2 s 120906 0 120962 800 6 la_data_out[96]
port 397 nsew signal output
rlabel metal2 s 121734 0 121790 800 6 la_data_out[97]
port 398 nsew signal output
rlabel metal2 s 122562 0 122618 800 6 la_data_out[98]
port 399 nsew signal output
rlabel metal2 s 123390 0 123446 800 6 la_data_out[99]
port 400 nsew signal output
rlabel metal2 s 48870 0 48926 800 6 la_data_out[9]
port 401 nsew signal output
rlabel metal2 s 41694 0 41750 800 6 la_oenb[0]
port 402 nsew signal input
rlabel metal2 s 124494 0 124550 800 6 la_oenb[100]
port 403 nsew signal input
rlabel metal2 s 125322 0 125378 800 6 la_oenb[101]
port 404 nsew signal input
rlabel metal2 s 126150 0 126206 800 6 la_oenb[102]
port 405 nsew signal input
rlabel metal2 s 126978 0 127034 800 6 la_oenb[103]
port 406 nsew signal input
rlabel metal2 s 127806 0 127862 800 6 la_oenb[104]
port 407 nsew signal input
rlabel metal2 s 128634 0 128690 800 6 la_oenb[105]
port 408 nsew signal input
rlabel metal2 s 129462 0 129518 800 6 la_oenb[106]
port 409 nsew signal input
rlabel metal2 s 130290 0 130346 800 6 la_oenb[107]
port 410 nsew signal input
rlabel metal2 s 131118 0 131174 800 6 la_oenb[108]
port 411 nsew signal input
rlabel metal2 s 131946 0 132002 800 6 la_oenb[109]
port 412 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 la_oenb[10]
port 413 nsew signal input
rlabel metal2 s 132774 0 132830 800 6 la_oenb[110]
port 414 nsew signal input
rlabel metal2 s 133602 0 133658 800 6 la_oenb[111]
port 415 nsew signal input
rlabel metal2 s 134430 0 134486 800 6 la_oenb[112]
port 416 nsew signal input
rlabel metal2 s 135258 0 135314 800 6 la_oenb[113]
port 417 nsew signal input
rlabel metal2 s 136086 0 136142 800 6 la_oenb[114]
port 418 nsew signal input
rlabel metal2 s 136914 0 136970 800 6 la_oenb[115]
port 419 nsew signal input
rlabel metal2 s 137742 0 137798 800 6 la_oenb[116]
port 420 nsew signal input
rlabel metal2 s 138570 0 138626 800 6 la_oenb[117]
port 421 nsew signal input
rlabel metal2 s 139398 0 139454 800 6 la_oenb[118]
port 422 nsew signal input
rlabel metal2 s 140226 0 140282 800 6 la_oenb[119]
port 423 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 la_oenb[11]
port 424 nsew signal input
rlabel metal2 s 141054 0 141110 800 6 la_oenb[120]
port 425 nsew signal input
rlabel metal2 s 141882 0 141938 800 6 la_oenb[121]
port 426 nsew signal input
rlabel metal2 s 142710 0 142766 800 6 la_oenb[122]
port 427 nsew signal input
rlabel metal2 s 143538 0 143594 800 6 la_oenb[123]
port 428 nsew signal input
rlabel metal2 s 144366 0 144422 800 6 la_oenb[124]
port 429 nsew signal input
rlabel metal2 s 145194 0 145250 800 6 la_oenb[125]
port 430 nsew signal input
rlabel metal2 s 146022 0 146078 800 6 la_oenb[126]
port 431 nsew signal input
rlabel metal2 s 146850 0 146906 800 6 la_oenb[127]
port 432 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 la_oenb[12]
port 433 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 la_oenb[13]
port 434 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 la_oenb[14]
port 435 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 la_oenb[15]
port 436 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 la_oenb[16]
port 437 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 la_oenb[17]
port 438 nsew signal input
rlabel metal2 s 56598 0 56654 800 6 la_oenb[18]
port 439 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 la_oenb[19]
port 440 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 la_oenb[1]
port 441 nsew signal input
rlabel metal2 s 58254 0 58310 800 6 la_oenb[20]
port 442 nsew signal input
rlabel metal2 s 59082 0 59138 800 6 la_oenb[21]
port 443 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 la_oenb[22]
port 444 nsew signal input
rlabel metal2 s 60738 0 60794 800 6 la_oenb[23]
port 445 nsew signal input
rlabel metal2 s 61566 0 61622 800 6 la_oenb[24]
port 446 nsew signal input
rlabel metal2 s 62394 0 62450 800 6 la_oenb[25]
port 447 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 la_oenb[26]
port 448 nsew signal input
rlabel metal2 s 64050 0 64106 800 6 la_oenb[27]
port 449 nsew signal input
rlabel metal2 s 64878 0 64934 800 6 la_oenb[28]
port 450 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 la_oenb[29]
port 451 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 la_oenb[2]
port 452 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 la_oenb[30]
port 453 nsew signal input
rlabel metal2 s 67362 0 67418 800 6 la_oenb[31]
port 454 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 la_oenb[32]
port 455 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 la_oenb[33]
port 456 nsew signal input
rlabel metal2 s 69846 0 69902 800 6 la_oenb[34]
port 457 nsew signal input
rlabel metal2 s 70674 0 70730 800 6 la_oenb[35]
port 458 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 la_oenb[36]
port 459 nsew signal input
rlabel metal2 s 72330 0 72386 800 6 la_oenb[37]
port 460 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 la_oenb[38]
port 461 nsew signal input
rlabel metal2 s 73986 0 74042 800 6 la_oenb[39]
port 462 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 la_oenb[3]
port 463 nsew signal input
rlabel metal2 s 74814 0 74870 800 6 la_oenb[40]
port 464 nsew signal input
rlabel metal2 s 75642 0 75698 800 6 la_oenb[41]
port 465 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 la_oenb[42]
port 466 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 la_oenb[43]
port 467 nsew signal input
rlabel metal2 s 78126 0 78182 800 6 la_oenb[44]
port 468 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 la_oenb[45]
port 469 nsew signal input
rlabel metal2 s 79782 0 79838 800 6 la_oenb[46]
port 470 nsew signal input
rlabel metal2 s 80610 0 80666 800 6 la_oenb[47]
port 471 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 la_oenb[48]
port 472 nsew signal input
rlabel metal2 s 82266 0 82322 800 6 la_oenb[49]
port 473 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 la_oenb[4]
port 474 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 la_oenb[50]
port 475 nsew signal input
rlabel metal2 s 83922 0 83978 800 6 la_oenb[51]
port 476 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 la_oenb[52]
port 477 nsew signal input
rlabel metal2 s 85578 0 85634 800 6 la_oenb[53]
port 478 nsew signal input
rlabel metal2 s 86406 0 86462 800 6 la_oenb[54]
port 479 nsew signal input
rlabel metal2 s 87234 0 87290 800 6 la_oenb[55]
port 480 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 la_oenb[56]
port 481 nsew signal input
rlabel metal2 s 88890 0 88946 800 6 la_oenb[57]
port 482 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_oenb[58]
port 483 nsew signal input
rlabel metal2 s 90546 0 90602 800 6 la_oenb[59]
port 484 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 la_oenb[5]
port 485 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 la_oenb[60]
port 486 nsew signal input
rlabel metal2 s 92202 0 92258 800 6 la_oenb[61]
port 487 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 la_oenb[62]
port 488 nsew signal input
rlabel metal2 s 93858 0 93914 800 6 la_oenb[63]
port 489 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 la_oenb[64]
port 490 nsew signal input
rlabel metal2 s 95514 0 95570 800 6 la_oenb[65]
port 491 nsew signal input
rlabel metal2 s 96342 0 96398 800 6 la_oenb[66]
port 492 nsew signal input
rlabel metal2 s 97170 0 97226 800 6 la_oenb[67]
port 493 nsew signal input
rlabel metal2 s 97998 0 98054 800 6 la_oenb[68]
port 494 nsew signal input
rlabel metal2 s 98826 0 98882 800 6 la_oenb[69]
port 495 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 la_oenb[6]
port 496 nsew signal input
rlabel metal2 s 99654 0 99710 800 6 la_oenb[70]
port 497 nsew signal input
rlabel metal2 s 100482 0 100538 800 6 la_oenb[71]
port 498 nsew signal input
rlabel metal2 s 101310 0 101366 800 6 la_oenb[72]
port 499 nsew signal input
rlabel metal2 s 102138 0 102194 800 6 la_oenb[73]
port 500 nsew signal input
rlabel metal2 s 102966 0 103022 800 6 la_oenb[74]
port 501 nsew signal input
rlabel metal2 s 103794 0 103850 800 6 la_oenb[75]
port 502 nsew signal input
rlabel metal2 s 104622 0 104678 800 6 la_oenb[76]
port 503 nsew signal input
rlabel metal2 s 105450 0 105506 800 6 la_oenb[77]
port 504 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 la_oenb[78]
port 505 nsew signal input
rlabel metal2 s 107106 0 107162 800 6 la_oenb[79]
port 506 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 la_oenb[7]
port 507 nsew signal input
rlabel metal2 s 107934 0 107990 800 6 la_oenb[80]
port 508 nsew signal input
rlabel metal2 s 108762 0 108818 800 6 la_oenb[81]
port 509 nsew signal input
rlabel metal2 s 109590 0 109646 800 6 la_oenb[82]
port 510 nsew signal input
rlabel metal2 s 110418 0 110474 800 6 la_oenb[83]
port 511 nsew signal input
rlabel metal2 s 111246 0 111302 800 6 la_oenb[84]
port 512 nsew signal input
rlabel metal2 s 112074 0 112130 800 6 la_oenb[85]
port 513 nsew signal input
rlabel metal2 s 112902 0 112958 800 6 la_oenb[86]
port 514 nsew signal input
rlabel metal2 s 113730 0 113786 800 6 la_oenb[87]
port 515 nsew signal input
rlabel metal2 s 114558 0 114614 800 6 la_oenb[88]
port 516 nsew signal input
rlabel metal2 s 115386 0 115442 800 6 la_oenb[89]
port 517 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 la_oenb[8]
port 518 nsew signal input
rlabel metal2 s 116214 0 116270 800 6 la_oenb[90]
port 519 nsew signal input
rlabel metal2 s 117042 0 117098 800 6 la_oenb[91]
port 520 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 la_oenb[92]
port 521 nsew signal input
rlabel metal2 s 118698 0 118754 800 6 la_oenb[93]
port 522 nsew signal input
rlabel metal2 s 119526 0 119582 800 6 la_oenb[94]
port 523 nsew signal input
rlabel metal2 s 120354 0 120410 800 6 la_oenb[95]
port 524 nsew signal input
rlabel metal2 s 121182 0 121238 800 6 la_oenb[96]
port 525 nsew signal input
rlabel metal2 s 122010 0 122066 800 6 la_oenb[97]
port 526 nsew signal input
rlabel metal2 s 122838 0 122894 800 6 la_oenb[98]
port 527 nsew signal input
rlabel metal2 s 123666 0 123722 800 6 la_oenb[99]
port 528 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 la_oenb[9]
port 529 nsew signal input
rlabel metal2 s 147126 0 147182 800 6 user_clock2
port 530 nsew signal input
rlabel metal2 s 147402 0 147458 800 6 user_irq[0]
port 531 nsew signal output
rlabel metal2 s 147678 0 147734 800 6 user_irq[1]
port 532 nsew signal output
rlabel metal2 s 147954 0 148010 800 6 user_irq[2]
port 533 nsew signal output
rlabel metal2 s 11886 0 11942 800 6 wb_clk_i
port 534 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 wb_rst_i
port 535 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wbs_ack_o
port 536 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 wbs_adr_i[0]
port 537 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 wbs_adr_i[10]
port 538 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 wbs_adr_i[11]
port 539 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 wbs_adr_i[12]
port 540 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 wbs_adr_i[13]
port 541 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 wbs_adr_i[14]
port 542 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 wbs_adr_i[15]
port 543 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 wbs_adr_i[16]
port 544 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 wbs_adr_i[17]
port 545 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 wbs_adr_i[18]
port 546 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 wbs_adr_i[19]
port 547 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 wbs_adr_i[1]
port 548 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 wbs_adr_i[20]
port 549 nsew signal input
rlabel metal2 s 32034 0 32090 800 6 wbs_adr_i[21]
port 550 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 wbs_adr_i[22]
port 551 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 wbs_adr_i[23]
port 552 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 wbs_adr_i[24]
port 553 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 wbs_adr_i[25]
port 554 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 wbs_adr_i[26]
port 555 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 wbs_adr_i[27]
port 556 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 wbs_adr_i[28]
port 557 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 wbs_adr_i[29]
port 558 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 wbs_adr_i[2]
port 559 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 wbs_adr_i[30]
port 560 nsew signal input
rlabel metal2 s 40314 0 40370 800 6 wbs_adr_i[31]
port 561 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 wbs_adr_i[3]
port 562 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_adr_i[4]
port 563 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 wbs_adr_i[5]
port 564 nsew signal input
rlabel metal2 s 19614 0 19670 800 6 wbs_adr_i[6]
port 565 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wbs_adr_i[7]
port 566 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 wbs_adr_i[8]
port 567 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 wbs_adr_i[9]
port 568 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 wbs_cyc_i
port 569 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_dat_i[0]
port 570 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 wbs_dat_i[10]
port 571 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 wbs_dat_i[11]
port 572 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 wbs_dat_i[12]
port 573 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 wbs_dat_i[13]
port 574 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 wbs_dat_i[14]
port 575 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 wbs_dat_i[15]
port 576 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 wbs_dat_i[16]
port 577 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 wbs_dat_i[17]
port 578 nsew signal input
rlabel metal2 s 29826 0 29882 800 6 wbs_dat_i[18]
port 579 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 wbs_dat_i[19]
port 580 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 wbs_dat_i[1]
port 581 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 wbs_dat_i[20]
port 582 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 wbs_dat_i[21]
port 583 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 wbs_dat_i[22]
port 584 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 wbs_dat_i[23]
port 585 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 wbs_dat_i[24]
port 586 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 wbs_dat_i[25]
port 587 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 wbs_dat_i[26]
port 588 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 wbs_dat_i[27]
port 589 nsew signal input
rlabel metal2 s 38106 0 38162 800 6 wbs_dat_i[28]
port 590 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 wbs_dat_i[29]
port 591 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 wbs_dat_i[2]
port 592 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 wbs_dat_i[30]
port 593 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 wbs_dat_i[31]
port 594 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 wbs_dat_i[3]
port 595 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 wbs_dat_i[4]
port 596 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 wbs_dat_i[5]
port 597 nsew signal input
rlabel metal2 s 19890 0 19946 800 6 wbs_dat_i[6]
port 598 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 wbs_dat_i[7]
port 599 nsew signal input
rlabel metal2 s 21546 0 21602 800 6 wbs_dat_i[8]
port 600 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 wbs_dat_i[9]
port 601 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 wbs_dat_o[0]
port 602 nsew signal output
rlabel metal2 s 23478 0 23534 800 6 wbs_dat_o[10]
port 603 nsew signal output
rlabel metal2 s 24306 0 24362 800 6 wbs_dat_o[11]
port 604 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 wbs_dat_o[12]
port 605 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 wbs_dat_o[13]
port 606 nsew signal output
rlabel metal2 s 26790 0 26846 800 6 wbs_dat_o[14]
port 607 nsew signal output
rlabel metal2 s 27618 0 27674 800 6 wbs_dat_o[15]
port 608 nsew signal output
rlabel metal2 s 28446 0 28502 800 6 wbs_dat_o[16]
port 609 nsew signal output
rlabel metal2 s 29274 0 29330 800 6 wbs_dat_o[17]
port 610 nsew signal output
rlabel metal2 s 30102 0 30158 800 6 wbs_dat_o[18]
port 611 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 wbs_dat_o[19]
port 612 nsew signal output
rlabel metal2 s 15198 0 15254 800 6 wbs_dat_o[1]
port 613 nsew signal output
rlabel metal2 s 31758 0 31814 800 6 wbs_dat_o[20]
port 614 nsew signal output
rlabel metal2 s 32586 0 32642 800 6 wbs_dat_o[21]
port 615 nsew signal output
rlabel metal2 s 33414 0 33470 800 6 wbs_dat_o[22]
port 616 nsew signal output
rlabel metal2 s 34242 0 34298 800 6 wbs_dat_o[23]
port 617 nsew signal output
rlabel metal2 s 35070 0 35126 800 6 wbs_dat_o[24]
port 618 nsew signal output
rlabel metal2 s 35898 0 35954 800 6 wbs_dat_o[25]
port 619 nsew signal output
rlabel metal2 s 36726 0 36782 800 6 wbs_dat_o[26]
port 620 nsew signal output
rlabel metal2 s 37554 0 37610 800 6 wbs_dat_o[27]
port 621 nsew signal output
rlabel metal2 s 38382 0 38438 800 6 wbs_dat_o[28]
port 622 nsew signal output
rlabel metal2 s 39210 0 39266 800 6 wbs_dat_o[29]
port 623 nsew signal output
rlabel metal2 s 16302 0 16358 800 6 wbs_dat_o[2]
port 624 nsew signal output
rlabel metal2 s 40038 0 40094 800 6 wbs_dat_o[30]
port 625 nsew signal output
rlabel metal2 s 40866 0 40922 800 6 wbs_dat_o[31]
port 626 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 wbs_dat_o[3]
port 627 nsew signal output
rlabel metal2 s 18510 0 18566 800 6 wbs_dat_o[4]
port 628 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 wbs_dat_o[5]
port 629 nsew signal output
rlabel metal2 s 20166 0 20222 800 6 wbs_dat_o[6]
port 630 nsew signal output
rlabel metal2 s 20994 0 21050 800 6 wbs_dat_o[7]
port 631 nsew signal output
rlabel metal2 s 21822 0 21878 800 6 wbs_dat_o[8]
port 632 nsew signal output
rlabel metal2 s 22650 0 22706 800 6 wbs_dat_o[9]
port 633 nsew signal output
rlabel metal2 s 14370 0 14426 800 6 wbs_sel_i[0]
port 634 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 wbs_sel_i[1]
port 635 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 wbs_sel_i[2]
port 636 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wbs_sel_i[3]
port 637 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 wbs_stb_i
port 638 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wbs_we_i
port 639 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 160000 160000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 16809442
string GDS_FILE /openlane/designs/fp_division/runs/RUN_2023.11.25_16.34.47/results/signoff/user_project_wrapper.magic.gds
string GDS_START 958998
<< end >>

