VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ks_vandana_fp_div
  CLASS BLOCK ;
  FOREIGN ks_vandana_fp_div ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 400.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 13.020 10.640 14.620 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.020 10.640 39.620 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 63.020 10.640 64.620 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.020 10.640 89.620 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 113.020 10.640 114.620 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.020 10.640 139.620 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 163.020 10.640 164.620 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.020 10.640 189.620 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 213.020 10.640 214.620 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 238.020 10.640 239.620 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 263.020 10.640 264.620 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 288.020 10.640 289.620 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 313.020 10.640 314.620 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 338.020 10.640 339.620 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 363.020 10.640 364.620 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 388.020 10.640 389.620 389.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 18.380 394.460 19.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 43.380 394.460 44.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 68.380 394.460 69.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 93.380 394.460 94.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 118.380 394.460 119.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 143.380 394.460 144.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 168.380 394.460 169.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 193.380 394.460 194.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 218.380 394.460 219.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 243.380 394.460 244.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 268.380 394.460 269.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 293.380 394.460 294.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 318.380 394.460 319.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 343.380 394.460 344.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 368.380 394.460 369.980 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.720 10.640 11.320 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 34.720 10.640 36.320 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 59.720 10.640 61.320 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 84.720 10.640 86.320 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 109.720 10.640 111.320 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 134.720 10.640 136.320 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 159.720 10.640 161.320 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.720 10.640 186.320 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 209.720 10.640 211.320 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 234.720 10.640 236.320 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 259.720 10.640 261.320 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 284.720 10.640 286.320 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 309.720 10.640 311.320 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.720 10.640 336.320 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 359.720 10.640 361.320 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 384.720 10.640 386.320 389.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 15.080 394.460 16.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 40.080 394.460 41.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 65.080 394.460 66.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 90.080 394.460 91.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 115.080 394.460 116.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 140.080 394.460 141.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 165.080 394.460 166.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 190.080 394.460 191.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 215.080 394.460 216.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 240.080 394.460 241.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 265.080 394.460 266.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 290.080 394.460 291.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 315.080 394.460 316.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 340.080 394.460 341.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 365.080 394.460 366.680 ;
    END
  END VPWR
  PIN a1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 396.000 167.810 399.000 ;
    END
  END a1[0]
  PIN a1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 396.000 248.310 399.000 ;
    END
  END a1[10]
  PIN a1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 272.040 4.000 272.640 ;
    END
  END a1[11]
  PIN a1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 391.040 4.000 391.640 ;
    END
  END a1[12]
  PIN a1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 1.000 322.370 4.000 ;
    END
  END a1[13]
  PIN a1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 1.000 96.970 4.000 ;
    END
  END a1[14]
  PIN a1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 396.000 151.710 399.000 ;
    END
  END a1[15]
  PIN a1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 238.040 4.000 238.640 ;
    END
  END a1[16]
  PIN a1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 187.040 4.000 187.640 ;
    END
  END a1[17]
  PIN a1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 1.000 48.670 4.000 ;
    END
  END a1[18]
  PIN a1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 0.040 399.000 0.640 ;
    END
  END a1[19]
  PIN a1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 306.040 399.000 306.640 ;
    END
  END a1[1]
  PIN a1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 1.000 370.670 4.000 ;
    END
  END a1[20]
  PIN a1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 396.000 393.210 399.000 ;
    END
  END a1[21]
  PIN a1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 170.040 399.000 170.640 ;
    END
  END a1[22]
  PIN a1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 1.000 145.270 4.000 ;
    END
  END a1[23]
  PIN a1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 357.040 399.000 357.640 ;
    END
  END a1[24]
  PIN a1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 396.000 119.510 399.000 ;
    END
  END a1[25]
  PIN a1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 323.040 399.000 323.640 ;
    END
  END a1[26]
  PIN a1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 374.040 399.000 374.640 ;
    END
  END a1[27]
  PIN a1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 1.000 225.770 4.000 ;
    END
  END a1[28]
  PIN a1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 396.000 280.510 399.000 ;
    END
  END a1[29]
  PIN a1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 204.040 399.000 204.640 ;
    END
  END a1[2]
  PIN a1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 102.040 399.000 102.640 ;
    END
  END a1[30]
  PIN a1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 51.040 4.000 51.640 ;
    END
  END a1[31]
  PIN a1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 1.000 161.370 4.000 ;
    END
  END a1[3]
  PIN a1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 1.000 338.470 4.000 ;
    END
  END a1[4]
  PIN a1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 396.000 183.910 399.000 ;
    END
  END a1[5]
  PIN a1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 396.000 264.410 399.000 ;
    END
  END a1[6]
  PIN a1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 340.040 399.000 340.640 ;
    END
  END a1[7]
  PIN a1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 68.040 399.000 68.640 ;
    END
  END a1[8]
  PIN a1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 396.000 200.010 399.000 ;
    END
  END a1[9]
  PIN b1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 396.000 6.810 399.000 ;
    END
  END b1[0]
  PIN b1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 396.000 344.910 399.000 ;
    END
  END b1[10]
  PIN b1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 1.000 80.870 4.000 ;
    END
  END b1[11]
  PIN b1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 396.000 135.610 399.000 ;
    END
  END b1[12]
  PIN b1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 289.040 399.000 289.640 ;
    END
  END b1[13]
  PIN b1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 119.040 399.000 119.640 ;
    END
  END b1[14]
  PIN b1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 396.000 232.210 399.000 ;
    END
  END b1[15]
  PIN b1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 396.000 361.010 399.000 ;
    END
  END b1[16]
  PIN b1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 1.000 386.770 4.000 ;
    END
  END b1[17]
  PIN b1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 272.040 399.000 272.640 ;
    END
  END b1[18]
  PIN b1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 289.040 4.000 289.640 ;
    END
  END b1[19]
  PIN b1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 1.000 257.970 4.000 ;
    END
  END b1[1]
  PIN b1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 204.040 4.000 204.640 ;
    END
  END b1[20]
  PIN b1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 51.040 399.000 51.640 ;
    END
  END b1[21]
  PIN b1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 17.040 4.000 17.640 ;
    END
  END b1[22]
  PIN b1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 374.040 4.000 374.640 ;
    END
  END b1[23]
  PIN b1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 323.040 4.000 323.640 ;
    END
  END b1[24]
  PIN b1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 306.040 4.000 306.640 ;
    END
  END b1[25]
  PIN b1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 1.000 290.170 4.000 ;
    END
  END b1[26]
  PIN b1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 340.040 4.000 340.640 ;
    END
  END b1[27]
  PIN b1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 396.000 55.110 399.000 ;
    END
  END b1[28]
  PIN b1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 1.000 32.570 4.000 ;
    END
  END b1[29]
  PIN b1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 1.000 113.070 4.000 ;
    END
  END b1[2]
  PIN b1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 1.000 354.570 4.000 ;
    END
  END b1[30]
  PIN b1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 153.040 399.000 153.640 ;
    END
  END b1[31]
  PIN b1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 85.040 399.000 85.640 ;
    END
  END b1[3]
  PIN b1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 68.040 4.000 68.640 ;
    END
  END b1[4]
  PIN b1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 34.040 4.000 34.640 ;
    END
  END b1[5]
  PIN b1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 17.040 399.000 17.640 ;
    END
  END b1[6]
  PIN b1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 396.000 71.210 399.000 ;
    END
  END b1[7]
  PIN b1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 136.040 399.000 136.640 ;
    END
  END b1[8]
  PIN b1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 170.040 4.000 170.640 ;
    END
  END b1[9]
  PIN c[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 1.000 306.270 4.000 ;
    END
  END c[0]
  PIN c[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 255.040 399.000 255.640 ;
    END
  END c[10]
  PIN c[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 85.040 4.000 85.640 ;
    END
  END c[11]
  PIN c[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 255.040 4.000 255.640 ;
    END
  END c[12]
  PIN c[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 1.000 193.570 4.000 ;
    END
  END c[13]
  PIN c[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 1.000 0.370 4.000 ;
    END
  END c[14]
  PIN c[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 1.000 241.870 4.000 ;
    END
  END c[15]
  PIN c[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 396.000 103.410 399.000 ;
    END
  END c[16]
  PIN c[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 396.000 216.110 399.000 ;
    END
  END c[17]
  PIN c[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 136.040 4.000 136.640 ;
    END
  END c[18]
  PIN c[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 396.000 22.910 399.000 ;
    END
  END c[19]
  PIN c[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 221.040 4.000 221.640 ;
    END
  END c[1]
  PIN c[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 1.000 16.470 4.000 ;
    END
  END c[20]
  PIN c[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 396.000 377.110 399.000 ;
    END
  END c[21]
  PIN c[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 396.000 296.610 399.000 ;
    END
  END c[22]
  PIN c[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 1.000 177.470 4.000 ;
    END
  END c[23]
  PIN c[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 391.040 399.000 391.640 ;
    END
  END c[24]
  PIN c[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 34.040 399.000 34.640 ;
    END
  END c[25]
  PIN c[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 102.040 4.000 102.640 ;
    END
  END c[26]
  PIN c[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 221.040 399.000 221.640 ;
    END
  END c[27]
  PIN c[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 1.000 64.770 4.000 ;
    END
  END c[28]
  PIN c[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 1.000 129.170 4.000 ;
    END
  END c[29]
  PIN c[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 153.040 4.000 153.640 ;
    END
  END c[2]
  PIN c[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 238.040 399.000 238.640 ;
    END
  END c[30]
  PIN c[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 1.000 209.670 4.000 ;
    END
  END c[31]
  PIN c[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 396.000 328.810 399.000 ;
    END
  END c[3]
  PIN c[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 396.000 312.710 399.000 ;
    END
  END c[4]
  PIN c[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 396.000 39.010 399.000 ;
    END
  END c[5]
  PIN c[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 396.000 87.310 399.000 ;
    END
  END c[6]
  PIN c[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 1.000 274.070 4.000 ;
    END
  END c[7]
  PIN c[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 119.040 4.000 119.640 ;
    END
  END c[8]
  PIN c[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 357.040 4.000 357.640 ;
    END
  END c[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 187.040 399.000 187.640 ;
    END
  END clk
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 394.220 389.045 ;
      LAYER met1 ;
        RECT 0.070 6.500 399.670 391.640 ;
      LAYER met2 ;
        RECT 0.100 395.720 6.250 396.170 ;
        RECT 7.090 395.720 22.350 396.170 ;
        RECT 23.190 395.720 38.450 396.170 ;
        RECT 39.290 395.720 54.550 396.170 ;
        RECT 55.390 395.720 70.650 396.170 ;
        RECT 71.490 395.720 86.750 396.170 ;
        RECT 87.590 395.720 102.850 396.170 ;
        RECT 103.690 395.720 118.950 396.170 ;
        RECT 119.790 395.720 135.050 396.170 ;
        RECT 135.890 395.720 151.150 396.170 ;
        RECT 151.990 395.720 167.250 396.170 ;
        RECT 168.090 395.720 183.350 396.170 ;
        RECT 184.190 395.720 199.450 396.170 ;
        RECT 200.290 395.720 215.550 396.170 ;
        RECT 216.390 395.720 231.650 396.170 ;
        RECT 232.490 395.720 247.750 396.170 ;
        RECT 248.590 395.720 263.850 396.170 ;
        RECT 264.690 395.720 279.950 396.170 ;
        RECT 280.790 395.720 296.050 396.170 ;
        RECT 296.890 395.720 312.150 396.170 ;
        RECT 312.990 395.720 328.250 396.170 ;
        RECT 329.090 395.720 344.350 396.170 ;
        RECT 345.190 395.720 360.450 396.170 ;
        RECT 361.290 395.720 376.550 396.170 ;
        RECT 377.390 395.720 392.650 396.170 ;
        RECT 393.490 395.720 399.650 396.170 ;
        RECT 0.100 4.280 399.650 395.720 ;
        RECT 0.650 0.720 15.910 4.280 ;
        RECT 16.750 0.720 32.010 4.280 ;
        RECT 32.850 0.720 48.110 4.280 ;
        RECT 48.950 0.720 64.210 4.280 ;
        RECT 65.050 0.720 80.310 4.280 ;
        RECT 81.150 0.720 96.410 4.280 ;
        RECT 97.250 0.720 112.510 4.280 ;
        RECT 113.350 0.720 128.610 4.280 ;
        RECT 129.450 0.720 144.710 4.280 ;
        RECT 145.550 0.720 160.810 4.280 ;
        RECT 161.650 0.720 176.910 4.280 ;
        RECT 177.750 0.720 193.010 4.280 ;
        RECT 193.850 0.720 209.110 4.280 ;
        RECT 209.950 0.720 225.210 4.280 ;
        RECT 226.050 0.720 241.310 4.280 ;
        RECT 242.150 0.720 257.410 4.280 ;
        RECT 258.250 0.720 273.510 4.280 ;
        RECT 274.350 0.720 289.610 4.280 ;
        RECT 290.450 0.720 305.710 4.280 ;
        RECT 306.550 0.720 321.810 4.280 ;
        RECT 322.650 0.720 337.910 4.280 ;
        RECT 338.750 0.720 354.010 4.280 ;
        RECT 354.850 0.720 370.110 4.280 ;
        RECT 370.950 0.720 386.210 4.280 ;
        RECT 387.050 0.720 399.650 4.280 ;
        RECT 0.100 0.155 399.650 0.720 ;
      LAYER met3 ;
        RECT 4.000 392.040 399.675 392.185 ;
        RECT 4.400 390.640 395.600 392.040 ;
        RECT 399.400 390.640 399.675 392.040 ;
        RECT 4.000 375.040 399.675 390.640 ;
        RECT 4.400 373.640 395.600 375.040 ;
        RECT 399.400 373.640 399.675 375.040 ;
        RECT 4.000 358.040 399.675 373.640 ;
        RECT 4.400 356.640 395.600 358.040 ;
        RECT 399.400 356.640 399.675 358.040 ;
        RECT 4.000 341.040 399.675 356.640 ;
        RECT 4.400 339.640 395.600 341.040 ;
        RECT 399.400 339.640 399.675 341.040 ;
        RECT 4.000 324.040 399.675 339.640 ;
        RECT 4.400 322.640 395.600 324.040 ;
        RECT 399.400 322.640 399.675 324.040 ;
        RECT 4.000 307.040 399.675 322.640 ;
        RECT 4.400 305.640 395.600 307.040 ;
        RECT 399.400 305.640 399.675 307.040 ;
        RECT 4.000 290.040 399.675 305.640 ;
        RECT 4.400 288.640 395.600 290.040 ;
        RECT 399.400 288.640 399.675 290.040 ;
        RECT 4.000 273.040 399.675 288.640 ;
        RECT 4.400 271.640 395.600 273.040 ;
        RECT 399.400 271.640 399.675 273.040 ;
        RECT 4.000 256.040 399.675 271.640 ;
        RECT 4.400 254.640 395.600 256.040 ;
        RECT 399.400 254.640 399.675 256.040 ;
        RECT 4.000 239.040 399.675 254.640 ;
        RECT 4.400 237.640 395.600 239.040 ;
        RECT 399.400 237.640 399.675 239.040 ;
        RECT 4.000 222.040 399.675 237.640 ;
        RECT 4.400 220.640 395.600 222.040 ;
        RECT 399.400 220.640 399.675 222.040 ;
        RECT 4.000 205.040 399.675 220.640 ;
        RECT 4.400 203.640 395.600 205.040 ;
        RECT 399.400 203.640 399.675 205.040 ;
        RECT 4.000 188.040 399.675 203.640 ;
        RECT 4.400 186.640 395.600 188.040 ;
        RECT 399.400 186.640 399.675 188.040 ;
        RECT 4.000 171.040 399.675 186.640 ;
        RECT 4.400 169.640 395.600 171.040 ;
        RECT 399.400 169.640 399.675 171.040 ;
        RECT 4.000 154.040 399.675 169.640 ;
        RECT 4.400 152.640 395.600 154.040 ;
        RECT 399.400 152.640 399.675 154.040 ;
        RECT 4.000 137.040 399.675 152.640 ;
        RECT 4.400 135.640 395.600 137.040 ;
        RECT 399.400 135.640 399.675 137.040 ;
        RECT 4.000 120.040 399.675 135.640 ;
        RECT 4.400 118.640 395.600 120.040 ;
        RECT 399.400 118.640 399.675 120.040 ;
        RECT 4.000 103.040 399.675 118.640 ;
        RECT 4.400 101.640 395.600 103.040 ;
        RECT 399.400 101.640 399.675 103.040 ;
        RECT 4.000 86.040 399.675 101.640 ;
        RECT 4.400 84.640 395.600 86.040 ;
        RECT 399.400 84.640 399.675 86.040 ;
        RECT 4.000 69.040 399.675 84.640 ;
        RECT 4.400 67.640 395.600 69.040 ;
        RECT 399.400 67.640 399.675 69.040 ;
        RECT 4.000 52.040 399.675 67.640 ;
        RECT 4.400 50.640 395.600 52.040 ;
        RECT 399.400 50.640 399.675 52.040 ;
        RECT 4.000 35.040 399.675 50.640 ;
        RECT 4.400 33.640 395.600 35.040 ;
        RECT 399.400 33.640 399.675 35.040 ;
        RECT 4.000 18.040 399.675 33.640 ;
        RECT 4.400 16.640 395.600 18.040 ;
        RECT 399.400 16.640 399.675 18.040 ;
        RECT 4.000 1.040 399.675 16.640 ;
        RECT 4.000 0.175 395.600 1.040 ;
        RECT 399.400 0.175 399.675 1.040 ;
      LAYER met4 ;
        RECT 41.695 389.600 377.825 392.185 ;
        RECT 41.695 10.240 59.320 389.600 ;
        RECT 61.720 10.240 62.620 389.600 ;
        RECT 65.020 10.240 84.320 389.600 ;
        RECT 86.720 10.240 87.620 389.600 ;
        RECT 90.020 10.240 109.320 389.600 ;
        RECT 111.720 10.240 112.620 389.600 ;
        RECT 115.020 10.240 134.320 389.600 ;
        RECT 136.720 10.240 137.620 389.600 ;
        RECT 140.020 10.240 159.320 389.600 ;
        RECT 161.720 10.240 162.620 389.600 ;
        RECT 165.020 10.240 184.320 389.600 ;
        RECT 186.720 10.240 187.620 389.600 ;
        RECT 190.020 10.240 209.320 389.600 ;
        RECT 211.720 10.240 212.620 389.600 ;
        RECT 215.020 10.240 234.320 389.600 ;
        RECT 236.720 10.240 237.620 389.600 ;
        RECT 240.020 10.240 259.320 389.600 ;
        RECT 261.720 10.240 262.620 389.600 ;
        RECT 265.020 10.240 284.320 389.600 ;
        RECT 286.720 10.240 287.620 389.600 ;
        RECT 290.020 10.240 309.320 389.600 ;
        RECT 311.720 10.240 312.620 389.600 ;
        RECT 315.020 10.240 334.320 389.600 ;
        RECT 336.720 10.240 337.620 389.600 ;
        RECT 340.020 10.240 359.320 389.600 ;
        RECT 361.720 10.240 362.620 389.600 ;
        RECT 365.020 10.240 377.825 389.600 ;
        RECT 41.695 7.655 377.825 10.240 ;
  END
END ks_vandana_fp_div
END LIBRARY

