* NGSPICE file created from user_project_wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_2 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4bb_2 abstract view
.subckt sky130_fd_sc_hd__nand4bb_2 A_N B_N C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_1 abstract view
.subckt sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_2 abstract view
.subckt sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

.subckt user_project_wrapper VGND VPWR analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[2]
+ analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7] analog_io[8] analog_io[9]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110]
+ la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115]
+ la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120]
+ la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125]
+ la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64]
+ la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75]
+ la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91]
+ la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97]
+ la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102]
+ la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109]
+ la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115]
+ la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121]
+ la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12]
+ la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19]
+ la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31]
+ la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38]
+ la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44]
+ la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50]
+ la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57]
+ la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63]
+ la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6]
+ la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76]
+ la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89]
+ la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95]
+ la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0]
+ user_irq[1] user_irq[2] wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
+ wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
+ wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4]
+ wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_246_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_268_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8235_ net66 net20 VGND VGND VPWR VPWR fd.a\[27\] sky130_fd_sc_hd__dfxtp_1
Xfd._5447_ fd._0518_ VGND VGND VPWR VPWR fd._0519_ sky130_fd_sc_hd__inv_2
XFILLER_210_1519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_269_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_255_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8166_ fd.a\[28\] fd._3480_ fd._3471_ VGND VGND VPWR VPWR fd._3481_ sky130_fd_sc_hd__a21oi_2
XFILLER_67_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5378_ fd._0125_ fd._0442_ VGND VGND VPWR VPWR fd._0443_ sky130_fd_sc_hd__nand2_1
XFILLER_270_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7117_ fd._2164_ VGND VGND VPWR VPWR fd._2356_ sky130_fd_sc_hd__clkinv_2
XFILLER_110_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4329_ fd._2738_ fd._2793_ VGND VGND VPWR VPWR fd._2804_ sky130_fd_sc_hd__nor2_1
XFILLER_208_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8097_ fd._0453_ fd._0651_ fd._3411_ VGND VGND VPWR VPWR fd._3418_ sky130_fd_sc_hd__mux2_1
XFILLER_39_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7048_ fd._0382_ fd._2098_ VGND VGND VPWR VPWR fd._2280_ sky130_fd_sc_hd__nor2_1
XFILLER_39_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_260_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_278_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4680_ fd._3592_ fd._3594_ fd._3599_ VGND VGND VPWR VPWR fd._3774_ sky130_fd_sc_hd__and3_1
XFILLER_194_1360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6350_ fd._1507_ fd._1510_ VGND VGND VPWR VPWR fd._1512_ sky130_fd_sc_hd__nor2_1
XFILLER_123_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_268_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5301_ fd._0292_ fd._0357_ VGND VGND VPWR VPWR fd._0358_ sky130_fd_sc_hd__nand2_1
XFILLER_284_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6281_ fd._1435_ fd._1292_ VGND VGND VPWR VPWR fd._1436_ sky130_fd_sc_hd__nand2_1
XFILLER_49_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_283_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._8020_ fd._3334_ fd._3199_ VGND VGND VPWR VPWR fd._3349_ sky130_fd_sc_hd__xnor2_1
XFILLER_64_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5232_ fd._0195_ fd._0281_ fd._0270_ VGND VGND VPWR VPWR fd._0282_ sky130_fd_sc_hd__mux2_1
XFILLER_168_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5163_ fd._0205_ VGND VGND VPWR VPWR fd._0206_ sky130_fd_sc_hd__inv_1
XFILLER_184_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4114_ fd.a\[7\] VGND VGND VPWR VPWR fd._0439_ sky130_fd_sc_hd__inv_2
XFILLER_166_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_1626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5094_ fd._0125_ fd._0128_ fd._0129_ fd._4011_ VGND VGND VPWR VPWR fd._0130_ sky130_fd_sc_hd__a211o_1
XFILLER_166_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7804_ fd._2093_ fd._3109_ VGND VGND VPWR VPWR fd._3111_ sky130_fd_sc_hd__nor2_1
XFILLER_285_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._5996_ fd._0952_ fd._1120_ fd._1046_ fd._1122_ VGND VGND VPWR VPWR fd._1123_ sky130_fd_sc_hd__a31oi_2
XFILLER_118_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_277_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4947_ fd._0846_ fd._4040_ VGND VGND VPWR VPWR fd._4041_ sky130_fd_sc_hd__nor2_1
XFILLER_173_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7735_ fd._2863_ fd._3033_ VGND VGND VPWR VPWR fd._3036_ sky130_fd_sc_hd__nand2_1
XFILLER_118_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7666_ fd._2763_ fd._2956_ fd._2959_ VGND VGND VPWR VPWR fd._2960_ sky130_fd_sc_hd__o21ba_1
XFILLER_271_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4878_ fd._1253_ fd._3971_ VGND VGND VPWR VPWR fd._3972_ sky130_fd_sc_hd__nand2_1
XFILLER_216_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6617_ fd._1802_ fd._1805_ fd._1637_ VGND VGND VPWR VPWR fd._1806_ sky130_fd_sc_hd__o21a_1
XFILLER_271_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7597_ fd._2880_ fd._2883_ fd._2877_ VGND VGND VPWR VPWR fd._2884_ sky130_fd_sc_hd__mux2_1
XFILLER_141_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6548_ fd._1722_ fd._1728_ VGND VGND VPWR VPWR fd._1730_ sky130_fd_sc_hd__and2_1
XFILLER_99_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6479_ fd._1453_ fd._1653_ fd._1615_ VGND VGND VPWR VPWR fd._1654_ sky130_fd_sc_hd__mux2_1
XFILLER_132_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8218_ net73 net2 VGND VGND VPWR VPWR fd.a\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_28_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8149_ fd._3450_ fd._3454_ fd._3462_ VGND VGND VPWR VPWR fd._3464_ sky130_fd_sc_hd__o21a_1
XFILLER_215_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_260_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_265_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5850_ fd._0724_ fd._0730_ VGND VGND VPWR VPWR fd._0962_ sky130_fd_sc_hd__xnor2_1
XFILLER_204_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_259_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4801_ fd._3708_ fd._3892_ VGND VGND VPWR VPWR fd._3895_ sky130_fd_sc_hd__nand2_1
XFILLER_183_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5781_ fd._0878_ fd._0884_ fd._0885_ VGND VGND VPWR VPWR fd._0886_ sky130_fd_sc_hd__o21a_1
XFILLER_154_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7520_ fd._1666_ fd._2702_ VGND VGND VPWR VPWR fd._2799_ sky130_fd_sc_hd__or2_1
XFILLER_115_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4732_ fd._3730_ fd._3788_ VGND VGND VPWR VPWR fd._3826_ sky130_fd_sc_hd__nand2_1
XFILLER_192_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7451_ fd._2720_ fd._2722_ VGND VGND VPWR VPWR fd._2723_ sky130_fd_sc_hd__xnor2_1
XFILLER_83_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4663_ fd._3628_ fd._3752_ fd._3756_ VGND VGND VPWR VPWR fd._3757_ sky130_fd_sc_hd__a21o_1
XFILLER_237_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6402_ fd._1390_ fd._1568_ VGND VGND VPWR VPWR fd._1569_ sky130_fd_sc_hd__and2_1
XFILLER_96_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7382_ fd._2447_ fd._2448_ fd._2444_ VGND VGND VPWR VPWR fd._2647_ sky130_fd_sc_hd__o21ai_1
XFILLER_29_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_257_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4594_ fd.b\[2\] VGND VGND VPWR VPWR fd._3688_ sky130_fd_sc_hd__buf_6
XFILLER_170_1639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_284_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6333_ fd._1482_ fd._1488_ fd._1491_ fd._1492_ VGND VGND VPWR VPWR fd._1493_ sky130_fd_sc_hd__a211o_1
XFILLER_211_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6264_ fd._1415_ fd._1416_ VGND VGND VPWR VPWR fd._1417_ sky130_fd_sc_hd__nor2_1
XFILLER_237_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8003_ fd._2566_ fd._3329_ VGND VGND VPWR VPWR fd._3330_ sky130_fd_sc_hd__and2_1
Xfd._5215_ fd._0240_ fd._0250_ fd._0262_ VGND VGND VPWR VPWR fd._0264_ sky130_fd_sc_hd__a21o_1
XFILLER_65_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6195_ fd._1318_ fd._1071_ fd._1052_ VGND VGND VPWR VPWR fd._1342_ sky130_fd_sc_hd__o21ai_1
XFILLER_20_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5146_ fd._1297_ fd._0187_ VGND VGND VPWR VPWR fd._0188_ sky130_fd_sc_hd__or2_1
XFILLER_212_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5077_ fd._0108_ fd._0111_ fd._0059_ VGND VGND VPWR VPWR fd._0112_ sky130_fd_sc_hd__mux2_2
XFILLER_221_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5979_ fd._1090_ fd._1096_ fd._1101_ fd._1103_ VGND VGND VPWR VPWR fd._1104_ sky130_fd_sc_hd__o31a_1
XFILLER_173_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7718_ fd._1685_ fd._3012_ VGND VGND VPWR VPWR fd._3017_ sky130_fd_sc_hd__or2_1
XFILLER_279_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7649_ fd._2937_ fd._2940_ fd._2874_ VGND VGND VPWR VPWR fd._2941_ sky130_fd_sc_hd__mux2_1
XFILLER_0_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_284_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_255_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_284_1236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_270_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_1704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_8599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_267_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5000_ fd._3808_ fd._3930_ VGND VGND VPWR VPWR fd._0027_ sky130_fd_sc_hd__or2_1
XFILLER_235_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_250_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_1590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_261_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_280_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._6951_ fd._2167_ fd._2172_ fd._2115_ VGND VGND VPWR VPWR fd._2173_ sky130_fd_sc_hd__mux2_1
XFILLER_261_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5902_ fd._0830_ fd._1018_ fd._0998_ VGND VGND VPWR VPWR fd._1019_ sky130_fd_sc_hd__mux2_1
XFILLER_187_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6882_ fd._1892_ fd._2096_ VGND VGND VPWR VPWR fd._2097_ sky130_fd_sc_hd__nor2_1
XFILLER_70_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5833_ fd._0707_ fd._0706_ VGND VGND VPWR VPWR fd._0943_ sky130_fd_sc_hd__nor2_1
XFILLER_200_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5764_ fd._0762_ fd._0866_ fd._0849_ VGND VGND VPWR VPWR fd._0867_ sky130_fd_sc_hd__mux2_1
XFILLER_192_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4715_ fd._3738_ fd._3741_ fd._3744_ VGND VGND VPWR VPWR fd._3809_ sky130_fd_sc_hd__a21o_1
Xfd._7503_ fd._2135_ fd._2776_ VGND VGND VPWR VPWR fd._2780_ sky130_fd_sc_hd__nor2_1
XFILLER_192_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5695_ fd._0789_ fd._0790_ VGND VGND VPWR VPWR fd._0792_ sky130_fd_sc_hd__nand2_1
XFILLER_157_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_272_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4646_ fd._3310_ fd._3739_ fd._3625_ VGND VGND VPWR VPWR fd._3740_ sky130_fd_sc_hd__mux2_1
XFILLER_170_1414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7434_ fd._2586_ fd._2593_ VGND VGND VPWR VPWR fd._2704_ sky130_fd_sc_hd__xnor2_1
XFILLER_269_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7365_ fd._1242_ fd._2627_ VGND VGND VPWR VPWR fd._2629_ sky130_fd_sc_hd__nand2_1
XFILLER_96_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4577_ fd._3668_ fd._3670_ VGND VGND VPWR VPWR fd._3671_ sky130_fd_sc_hd__nand2_1
XFILLER_57_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_284_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6316_ fd._1118_ fd._1474_ VGND VGND VPWR VPWR fd._1475_ sky130_fd_sc_hd__nor2_1
XFILLER_111_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7296_ fd._1211_ fd._1764_ fd._2423_ VGND VGND VPWR VPWR fd._2553_ sky130_fd_sc_hd__or3_1
XFILLER_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6247_ fd._0437_ fd._1340_ fd._1348_ VGND VGND VPWR VPWR fd._1399_ sky130_fd_sc_hd__and3_1
XFILLER_253_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_1529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_252_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_253_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6178_ fd._1322_ VGND VGND VPWR VPWR fd._1323_ sky130_fd_sc_hd__inv_2
XFILLER_240_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5129_ fd._4042_ fd._4046_ VGND VGND VPWR VPWR fd._0169_ sky130_fd_sc_hd__nand2_1
XFILLER_12_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_257_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_276_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_251_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_262_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_9086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_1518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4500_ fd._3565_ fd._3575_ fd._3583_ fd._3593_ VGND VGND VPWR VPWR fd._3594_ sky130_fd_sc_hd__nand4_1
XTAP_8396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5480_ fd._0550_ fd._3833_ fd._0554_ VGND VGND VPWR VPWR fd._0555_ sky130_fd_sc_hd__mux2_1
XFILLER_285_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_267_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4431_ fd._1979_ fd._3524_ VGND VGND VPWR VPWR fd._3525_ sky130_fd_sc_hd__nand2_1
XTAP_6961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7150_ fd._2149_ fd._2391_ fd._2322_ VGND VGND VPWR VPWR fd._2392_ sky130_fd_sc_hd__mux2_1
XFILLER_282_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4362_ fd.a\[22\] fd.b\[22\] VGND VGND VPWR VPWR fd._3167_ sky130_fd_sc_hd__and2_1
XFILLER_130_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6101_ fd._1126_ fd._1125_ VGND VGND VPWR VPWR fd._1238_ sky130_fd_sc_hd__or2_1
XFILLER_281_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7081_ fd._2315_ fd._2245_ VGND VGND VPWR VPWR fd._2316_ sky130_fd_sc_hd__nor2_1
Xfd._4293_ fd._1528_ fd._2375_ fd._2397_ VGND VGND VPWR VPWR fd._2408_ sky130_fd_sc_hd__a21oi_1
XFILLER_235_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6032_ fd._0482_ fd._1161_ VGND VGND VPWR VPWR fd._1162_ sky130_fd_sc_hd__nand2_1
XFILLER_130_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_1426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7983_ fd._3306_ fd._3292_ fd._3305_ fd._3303_ fd._3304_ VGND VGND VPWR VPWR fd._3308_
+ sky130_fd_sc_hd__o32a_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6934_ fd._1983_ fd._2143_ VGND VGND VPWR VPWR fd._2154_ sky130_fd_sc_hd__and2_1
XFILLER_147_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6865_ fd._1879_ fd._1884_ fd._2077_ VGND VGND VPWR VPWR fd._2079_ sky130_fd_sc_hd__a21oi_1
XFILLER_163_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5816_ fd._0526_ fd._0924_ VGND VGND VPWR VPWR fd._0925_ sky130_fd_sc_hd__nor2_1
XFILLER_115_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6796_ fd._0343_ fd._2002_ VGND VGND VPWR VPWR fd._2003_ sky130_fd_sc_hd__nand2_1
XFILLER_116_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5747_ fd._0848_ VGND VGND VPWR VPWR fd._0849_ sky130_fd_sc_hd__buf_6
XFILLER_217_1620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_258_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5678_ fd._0772_ fd._0608_ VGND VGND VPWR VPWR fd._0773_ sky130_fd_sc_hd__xnor2_1
XFILLER_135_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_269_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4629_ fd._3651_ fd._3715_ fd._3721_ fd._3722_ VGND VGND VPWR VPWR fd._3723_ sky130_fd_sc_hd__o31ai_1
Xfd._7417_ fd._2685_ fd._2614_ VGND VGND VPWR VPWR fd._2686_ sky130_fd_sc_hd__xnor2_1
XFILLER_285_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_285_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_268_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7348_ fd._2412_ fd._2609_ VGND VGND VPWR VPWR fd._2610_ sky130_fd_sc_hd__xnor2_1
XTAP_3609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_284_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7279_ fd._2384_ fd._2367_ VGND VGND VPWR VPWR fd._2534_ sky130_fd_sc_hd__or2b_1
XFILLER_26_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_272_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_285_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_1613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_279_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_283_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_264_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_263_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_268_1551 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_1584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._4980_ fd._2584_ fd._0003_ VGND VGND VPWR VPWR fd._0005_ sky130_fd_sc_hd__and2_1
XPHY_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_5 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfd._6650_ fd._1304_ fd._1841_ VGND VGND VPWR VPWR fd._1842_ sky130_fd_sc_hd__nor2_1
XFILLER_67_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5601_ fd._0683_ fd._0684_ fd._0685_ fd._0686_ fd._0687_ VGND VGND VPWR VPWR fd._0688_
+ sky130_fd_sc_hd__a311o_1
XFILLER_193_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6581_ fd._1626_ fd._1644_ fd._1718_ fd._1765_ fd._1590_ VGND VGND VPWR VPWR fd._1766_
+ sky130_fd_sc_hd__a32o_1
XTAP_8160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5532_ fd._0601_ fd._0606_ fd._0611_ fd._0478_ fd._0454_ VGND VGND VPWR VPWR fd._0612_
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_125_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1662 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8251_ net73 net3 VGND VGND VPWR VPWR fd.b\[11\] sky130_fd_sc_hd__dfxtp_2
Xfd._5463_ fd._0501_ fd._0535_ VGND VGND VPWR VPWR fd._0536_ sky130_fd_sc_hd__and2_1
XFILLER_6_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4414_ fd.b\[6\] fd._3507_ VGND VGND VPWR VPWR fd._3508_ sky130_fd_sc_hd__or2_1
XFILLER_227_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7202_ fd._2438_ VGND VGND VPWR VPWR fd._2449_ sky130_fd_sc_hd__inv_2
XFILLER_132_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_267_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8182_ net77 fd.mc\[6\] VGND VGND VPWR VPWR fd.c\[6\] sky130_fd_sc_hd__dfxtp_1
Xfd._5394_ fd._3947_ fd._0459_ VGND VGND VPWR VPWR fd._0460_ sky130_fd_sc_hd__or2_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_266_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7133_ fd._2368_ fd._2372_ fd._2322_ VGND VGND VPWR VPWR fd._2373_ sky130_fd_sc_hd__mux2_1
Xfd._4345_ fd.b\[18\] fd._2947_ VGND VGND VPWR VPWR fd._2980_ sky130_fd_sc_hd__xnor2_1
XFILLER_254_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_212_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_282_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7064_ fd._2291_ fd._2295_ fd._2296_ VGND VGND VPWR VPWR fd._2297_ sky130_fd_sc_hd__a21oi_2
XFILLER_81_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4276_ fd._2199_ fd._2210_ VGND VGND VPWR VPWR fd._2221_ sky130_fd_sc_hd__or2_1
XFILLER_207_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_project_wrapper_81 VGND VGND VPWR VPWR user_project_wrapper_81/HI io_oeb[3]
+ sky130_fd_sc_hd__conb_1
XFILLER_78_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_92 VGND VGND VPWR VPWR user_project_wrapper_92/HI io_oeb[14]
+ sky130_fd_sc_hd__conb_1
Xfd._6015_ fd._0968_ fd._1142_ VGND VGND VPWR VPWR fd._1144_ sky130_fd_sc_hd__nand2_1
XFILLER_35_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7966_ fd._3175_ fd._3289_ VGND VGND VPWR VPWR fd._3290_ sky130_fd_sc_hd__or2_1
XFILLER_202_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6917_ fd._1940_ VGND VGND VPWR VPWR fd._2136_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_148_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7897_ fd._3080_ fd._3213_ VGND VGND VPWR VPWR fd._3214_ sky130_fd_sc_hd__nand2_1
XFILLER_11_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6848_ fd._2057_ fd._2059_ VGND VGND VPWR VPWR fd._2060_ sky130_fd_sc_hd__xnor2_1
XFILLER_163_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6779_ fd._1559_ fd._1947_ VGND VGND VPWR VPWR fd._1984_ sky130_fd_sc_hd__or2_1
XFILLER_143_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_277_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_277_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_project_wrapper_108 VGND VGND VPWR VPWR user_project_wrapper_108/HI io_oeb[30]
+ sky130_fd_sc_hd__conb_1
XFILLER_33_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_119 VGND VGND VPWR VPWR user_project_wrapper_119/HI io_out[35]
+ sky130_fd_sc_hd__conb_1
XFILLER_120_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_218_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput42 net42 VGND VGND VPWR VPWR io_out[17] sky130_fd_sc_hd__buf_2
XFILLER_68_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput53 net53 VGND VGND VPWR VPWR io_out[27] sky130_fd_sc_hd__buf_2
XFILLER_194_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput64 net64 VGND VGND VPWR VPWR io_out[8] sky130_fd_sc_hd__buf_2
XFILLER_122_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_270_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4130_ fd.a\[8\] fd.b\[8\] VGND VGND VPWR VPWR fd._0615_ sky130_fd_sc_hd__nor2b_1
XFILLER_251_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_264_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_251_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7820_ fd._2973_ fd._2971_ VGND VGND VPWR VPWR fd._3129_ sky130_fd_sc_hd__and2b_1
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_1576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7751_ fd._3022_ VGND VGND VPWR VPWR fd._3053_ sky130_fd_sc_hd__inv_2
XFILLER_258_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4963_ fd._3831_ fd._3960_ VGND VGND VPWR VPWR fd._4058_ sky130_fd_sc_hd__nor2_1
XFILLER_172_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6702_ fd._1897_ fd._1856_ VGND VGND VPWR VPWR fd._1899_ sky130_fd_sc_hd__nor2b_1
XFILLER_51_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4894_ fd._3669_ fd._3987_ VGND VGND VPWR VPWR fd._3988_ sky130_fd_sc_hd__or2_1
XFILLER_172_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7682_ fd._2908_ fd._2920_ fd._2976_ fd._2906_ VGND VGND VPWR VPWR fd._2977_ sky130_fd_sc_hd__a31o_1
XFILLER_274_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6633_ fd._1636_ fd._1822_ fd._1813_ VGND VGND VPWR VPWR fd._1823_ sky130_fd_sc_hd__mux2_1
XFILLER_132_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6564_ fd._1575_ fd._1593_ VGND VGND VPWR VPWR fd._1747_ sky130_fd_sc_hd__xnor2_1
XFILLER_119_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_259_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5515_ fd._3580_ VGND VGND VPWR VPWR fd._0594_ sky130_fd_sc_hd__buf_6
XFILLER_268_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6495_ fd._1474_ fd._1670_ fd._1615_ VGND VGND VPWR VPWR fd._1672_ sky130_fd_sc_hd__mux2_1
XFILLER_119_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_269_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8234_ net66 net19 VGND VGND VPWR VPWR fd.a\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_234_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5446_ fd._0323_ fd._0517_ fd._0425_ VGND VGND VPWR VPWR fd._0518_ sky130_fd_sc_hd__mux2_1
XFILLER_214_1678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_283_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_269_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5377_ fd._0438_ fd._0441_ fd._0425_ VGND VGND VPWR VPWR fd._0442_ sky130_fd_sc_hd__mux2_1
Xfd._8165_ fd.b\[28\] VGND VGND VPWR VPWR fd._3480_ sky130_fd_sc_hd__inv_2
XFILLER_55_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4328_ fd.a\[21\] fd._2782_ fd._1231_ VGND VGND VPWR VPWR fd._2793_ sky130_fd_sc_hd__mux2_1
XFILLER_243_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7116_ fd._0504_ fd._2354_ VGND VGND VPWR VPWR fd._2355_ sky130_fd_sc_hd__nand2_1
XFILLER_247_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8096_ fd._3417_ VGND VGND VPWR VPWR fd.mc\[15\] sky130_fd_sc_hd__clkbuf_1
XFILLER_247_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_270_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4259_ fd._0252_ fd._1748_ VGND VGND VPWR VPWR fd._2034_ sky130_fd_sc_hd__nor2_1
XFILLER_223_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7047_ fd._2083_ fd._2095_ VGND VGND VPWR VPWR fd._2279_ sky130_fd_sc_hd__nor2_1
XFILLER_35_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_280_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7949_ fd._0821_ fd._3268_ VGND VGND VPWR VPWR fd._3271_ sky130_fd_sc_hd__or2_1
XFILLER_109_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_277_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_259_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5300_ fd._3833_ fd._0291_ VGND VGND VPWR VPWR fd._0357_ sky130_fd_sc_hd__nand2_1
XFILLER_7_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6280_ fd._1241_ fd._1283_ fd._1289_ fd._1293_ VGND VGND VPWR VPWR fd._1435_ sky130_fd_sc_hd__a31o_1
XTAP_5150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5231_ fd._0967_ fd._0196_ VGND VGND VPWR VPWR fd._0281_ sky130_fd_sc_hd__xnor2_1
XFILLER_209_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5162_ fd._0204_ fd._3971_ fd._0067_ VGND VGND VPWR VPWR fd._0205_ sky130_fd_sc_hd__mux2_1
XTAP_4493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4113_ fd.b\[7\] VGND VGND VPWR VPWR fd._0428_ sky130_fd_sc_hd__buf_2
XFILLER_75_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5093_ fd._3689_ fd._0050_ fd._0052_ fd._0057_ VGND VGND VPWR VPWR fd._0129_ sky130_fd_sc_hd__and4_1
XFILLER_17_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7803_ fd._2093_ fd._3109_ VGND VGND VPWR VPWR fd._3110_ sky130_fd_sc_hd__and2_1
XFILLER_242_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5995_ fd._0902_ fd._1046_ VGND VGND VPWR VPWR fd._1122_ sky130_fd_sc_hd__nor2_1
XFILLER_157_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7734_ fd._2863_ fd._3033_ VGND VGND VPWR VPWR fd._3034_ sky130_fd_sc_hd__or2_1
XFILLER_121_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4946_ fd._4038_ VGND VGND VPWR VPWR fd._4040_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_12_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7665_ fd._1764_ fd._2874_ fd._1211_ VGND VGND VPWR VPWR fd._2959_ sky130_fd_sc_hd__o21a_1
XFILLER_133_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4877_ fd._3816_ fd._3970_ fd._3961_ VGND VGND VPWR VPWR fd._3971_ sky130_fd_sc_hd__mux2_1
XFILLER_173_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6616_ fd._1804_ VGND VGND VPWR VPWR fd._1805_ sky130_fd_sc_hd__inv_2
XFILLER_173_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7596_ fd._2821_ fd._2882_ VGND VGND VPWR VPWR fd._2883_ sky130_fd_sc_hd__nand2_1
XFILLER_86_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6547_ fd._1722_ fd._1728_ VGND VGND VPWR VPWR fd._1729_ sky130_fd_sc_hd__nor2_1
XFILLER_134_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6478_ fd._1652_ VGND VGND VPWR VPWR fd._1653_ sky130_fd_sc_hd__inv_2
XFILLER_210_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8217_ net73 net32 VGND VGND VPWR VPWR fd.a\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_255_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5429_ fd._0330_ fd._0498_ VGND VGND VPWR VPWR fd._0499_ sky130_fd_sc_hd__xnor2_1
XFILLER_67_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_283_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8148_ fd._3450_ fd._3454_ fd._3462_ VGND VGND VPWR VPWR fd._3463_ sky130_fd_sc_hd__nor3_1
XFILLER_250_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8079_ fd._3406_ VGND VGND VPWR VPWR fd.mc\[7\] sky130_fd_sc_hd__clkbuf_1
XFILLER_36_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_282_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_259_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_1523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_278_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_1355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4800_ fd._3852_ fd._3846_ VGND VGND VPWR VPWR fd._3894_ sky130_fd_sc_hd__nor2_1
Xfd._5780_ fd._0482_ fd._0877_ VGND VGND VPWR VPWR fd._0885_ sky130_fd_sc_hd__nand2_1
XFILLER_10_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4731_ fd._3728_ fd._3824_ VGND VGND VPWR VPWR fd._3825_ sky130_fd_sc_hd__xnor2_1
XFILLER_170_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7450_ fd._2523_ fd._2721_ VGND VGND VPWR VPWR fd._2722_ sky130_fd_sc_hd__nand2_1
Xfd._4662_ fd._3035_ fd._3755_ VGND VGND VPWR VPWR fd._3756_ sky130_fd_sc_hd__xnor2_1
XFILLER_135_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._6401_ fd._0318_ fd._1391_ VGND VGND VPWR VPWR fd._1568_ sky130_fd_sc_hd__nand2_1
XFILLER_123_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4593_ fd.b\[3\] fd._3686_ VGND VGND VPWR VPWR fd._3687_ sky130_fd_sc_hd__nand2_1
XFILLER_155_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7381_ fd._2055_ fd._2616_ fd._2621_ VGND VGND VPWR VPWR fd._2646_ sky130_fd_sc_hd__mux2_1
XFILLER_25_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6332_ fd._1319_ fd._1487_ VGND VGND VPWR VPWR fd._1492_ sky130_fd_sc_hd__nor2_1
XFILLER_96_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_284_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6263_ fd._0916_ fd._1350_ VGND VGND VPWR VPWR fd._1416_ sky130_fd_sc_hd__nor2_1
XFILLER_49_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8002_ fd._3131_ fd._3328_ fd._3240_ VGND VGND VPWR VPWR fd._3329_ sky130_fd_sc_hd__mux2_1
XFILLER_20_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5214_ fd._3869_ VGND VGND VPWR VPWR fd._0262_ sky130_fd_sc_hd__buf_6
XFILLER_253_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6194_ fd._1303_ fd._1307_ fd._1323_ fd._1337_ fd._1339_ VGND VGND VPWR VPWR fd._1340_
+ sky130_fd_sc_hd__o2111ai_4
XTAP_4290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5145_ fd._0183_ fd._0184_ fd._0067_ fd._0185_ VGND VGND VPWR VPWR fd._0187_ sky130_fd_sc_hd__o31a_1
XFILLER_253_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_252_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5076_ fd._0110_ VGND VGND VPWR VPWR fd._0111_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_178_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_277_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5978_ fd._1102_ fd._1100_ VGND VGND VPWR VPWR fd._1103_ sky130_fd_sc_hd__nand2_1
XFILLER_134_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7717_ fd._1494_ fd._2891_ VGND VGND VPWR VPWR fd._3016_ sky130_fd_sc_hd__or2_1
XFILLER_273_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4929_ fd._3857_ fd._4022_ fd._3959_ VGND VGND VPWR VPWR fd._4023_ sky130_fd_sc_hd__mux2_1
XFILLER_118_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._7648_ fd._2938_ fd._2939_ VGND VGND VPWR VPWR fd._2940_ sky130_fd_sc_hd__xnor2_1
XTAP_6609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_project_wrapper_280 VGND VGND VPWR VPWR user_project_wrapper_280/HI wbs_dat_o[26]
+ sky130_fd_sc_hd__conb_1
XFILLER_47_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7579_ fd._2863_ fd._2861_ VGND VGND VPWR VPWR fd._2864_ sky130_fd_sc_hd__nor2_1
XFILLER_275_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_260_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_9202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_9213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_254_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_281_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_219_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_267_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_261_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._6950_ fd._2170_ fd._2171_ VGND VGND VPWR VPWR fd._2172_ sky130_fd_sc_hd__or2_1
XFILLER_128_1586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_261_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5901_ fd._0832_ fd._1017_ VGND VGND VPWR VPWR fd._1018_ sky130_fd_sc_hd__xnor2_1
XFILLER_175_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6881_ fd._1871_ fd._1886_ fd._1890_ VGND VGND VPWR VPWR fd._2096_ sky130_fd_sc_hd__and3_1
XFILLER_204_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5832_ fd._0918_ fd._0935_ fd._0940_ fd._0941_ VGND VGND VPWR VPWR fd._0942_ sky130_fd_sc_hd__a31o_1
XFILLER_204_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5763_ fd._0864_ fd._0865_ VGND VGND VPWR VPWR fd._0866_ sky130_fd_sc_hd__xor2_1
XFILLER_171_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7502_ fd._2726_ fd._2718_ VGND VGND VPWR VPWR fd._2779_ sky130_fd_sc_hd__and2b_1
XFILLER_83_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4714_ fd._3580_ fd._3807_ VGND VGND VPWR VPWR fd._3808_ sky130_fd_sc_hd__and2_1
XFILLER_196_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5694_ fd._3947_ fd._0788_ VGND VGND VPWR VPWR fd._0790_ sky130_fd_sc_hd__or2_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_272_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7433_ fd._1666_ fd._2702_ VGND VGND VPWR VPWR fd._2703_ sky130_fd_sc_hd__nand2_1
Xfd._4645_ fd._3449_ fd._3641_ VGND VGND VPWR VPWR fd._3739_ sky130_fd_sc_hd__xor2_1
XFILLER_142_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_272_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7364_ fd._2486_ fd._2623_ fd._2626_ VGND VGND VPWR VPWR fd._2627_ sky130_fd_sc_hd__o21a_1
XFILLER_97_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_284_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4576_ fd._3669_ fd._3667_ VGND VGND VPWR VPWR fd._3670_ sky130_fd_sc_hd__nand2_1
XFILLER_211_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6315_ fd._1245_ fd._1472_ fd._1422_ VGND VGND VPWR VPWR fd._1474_ sky130_fd_sc_hd__mux2_1
XFILLER_250_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_284_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7295_ fd._0318_ fd._2550_ VGND VGND VPWR VPWR fd._2552_ sky130_fd_sc_hd__or2_1
XFILLER_226_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6246_ fd._1393_ fd._1395_ fd._1397_ VGND VGND VPWR VPWR fd._1398_ sky130_fd_sc_hd__o21ai_1
XFILLER_42_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_253_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6177_ fd._1316_ fd._1321_ VGND VGND VPWR VPWR fd._1322_ sky130_fd_sc_hd__or2_1
XFILLER_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_253_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._5128_ fd._3833_ fd._0166_ fd._0167_ VGND VGND VPWR VPWR fd._0168_ sky130_fd_sc_hd__a21o_1
XFILLER_209_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_283_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5059_ fd._3999_ fd._4015_ VGND VGND VPWR VPWR fd._0092_ sky130_fd_sc_hd__or2_1
XFILLER_209_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_256_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_251_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_251_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_263_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_245_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_262_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_223_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_1647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1494 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_9087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4430_ fd.b\[1\] fd._3523_ VGND VGND VPWR VPWR fd._3524_ sky130_fd_sc_hd__nand2_1
XTAP_6962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_266_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4361_ fd._2804_ fd._3134_ fd._3145_ VGND VGND VPWR VPWR fd._3156_ sky130_fd_sc_hd__o21ai_1
XFILLER_130_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_266_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6100_ fd._0965_ fd._1236_ VGND VGND VPWR VPWR fd._1237_ sky130_fd_sc_hd__or2_1
XFILLER_47_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._4292_ fd._1440_ fd._2386_ VGND VGND VPWR VPWR fd._2397_ sky130_fd_sc_hd__or2_1
Xfd._7080_ fd._1816_ fd._2244_ VGND VGND VPWR VPWR fd._2315_ sky130_fd_sc_hd__and2_1
XFILLER_219_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6031_ fd._0594_ fd._1156_ fd._1160_ VGND VGND VPWR VPWR fd._1161_ sky130_fd_sc_hd__mux2_1
XFILLER_250_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_267_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_280_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_280_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._7982_ fd._3281_ fd._3293_ fd._3305_ fd._3306_ VGND VGND VPWR VPWR fd._3307_ sky130_fd_sc_hd__or4b_1
XFILLER_124_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_1438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6933_ fd._1955_ VGND VGND VPWR VPWR fd._2153_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_148_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6864_ fd._1871_ fd._1885_ VGND VGND VPWR VPWR fd._2077_ sky130_fd_sc_hd__nand2_1
XFILLER_141_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5815_ fd._0922_ VGND VGND VPWR VPWR fd._0924_ sky130_fd_sc_hd__inv_2
XFILLER_116_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._6795_ fd._1782_ fd._1969_ fd._2000_ VGND VGND VPWR VPWR fd._2002_ sky130_fd_sc_hd__a21oi_1
XFILLER_196_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_1367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5746_ fd._0801_ VGND VGND VPWR VPWR fd._0848_ sky130_fd_sc_hd__buf_6
XFILLER_157_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_277_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5677_ fd._0601_ fd._0606_ VGND VGND VPWR VPWR fd._0772_ sky130_fd_sc_hd__nor2_1
XFILLER_174_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7416_ fd._2615_ fd._2509_ VGND VGND VPWR VPWR fd._2685_ sky130_fd_sc_hd__or2b_1
Xfd._4628_ fd._3716_ fd._3720_ VGND VGND VPWR VPWR fd._3722_ sky130_fd_sc_hd__nand2_1
XFILLER_58_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_1529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_269_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7347_ fd._2417_ fd._2416_ VGND VGND VPWR VPWR fd._2609_ sky130_fd_sc_hd__or2b_1
XFILLER_135_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._4559_ fd._3495_ fd._3652_ fd._3625_ VGND VGND VPWR VPWR fd._3653_ sky130_fd_sc_hd__mux2_1
XFILLER_245_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7278_ fd._1559_ VGND VGND VPWR VPWR fd._2533_ sky130_fd_sc_hd__buf_6
XFILLER_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6229_ fd._0318_ fd._1204_ VGND VGND VPWR VPWR fd._1379_ sky130_fd_sc_hd__nand2_1
XFILLER_168_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_244_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_257_1467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1634 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_270_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_264_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_1530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_1503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_1558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_262_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_6 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5600_ fd._1341_ fd._0680_ VGND VGND VPWR VPWR fd._0687_ sky130_fd_sc_hd__and2_1
XFILLER_275_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._6580_ fd._1211_ fd._1764_ fd._1617_ VGND VGND VPWR VPWR fd._1765_ sky130_fd_sc_hd__or3_1
XFILLER_271_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_259_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5531_ fd._0608_ fd._0610_ VGND VGND VPWR VPWR fd._0611_ sky130_fd_sc_hd__nor2_1
XFILLER_3_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8250_ net73 net2 VGND VGND VPWR VPWR fd.b\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_234_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5462_ fd._3980_ fd._0500_ VGND VGND VPWR VPWR fd._0535_ sky130_fd_sc_hd__nand2_1
XFILLER_136_1674 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7201_ fd._2076_ fd._2418_ fd._2325_ VGND VGND VPWR VPWR fd._2448_ sky130_fd_sc_hd__mux2_1
XFILLER_121_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4413_ fd._1737_ fd._3506_ fd._3200_ VGND VGND VPWR VPWR fd._3507_ sky130_fd_sc_hd__mux2_1
XFILLER_234_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._8181_ net77 fd.mc\[5\] VGND VGND VPWR VPWR fd.c\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_94_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5393_ fd._0415_ fd._0458_ fd._0453_ VGND VGND VPWR VPWR fd._0459_ sky130_fd_sc_hd__mux2_1
XFILLER_39_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7132_ fd._2369_ fd._2371_ VGND VGND VPWR VPWR fd._2372_ sky130_fd_sc_hd__xnor2_1
XFILLER_43_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4344_ fd.b\[18\] fd._2925_ fd._2947_ fd._2958_ VGND VGND VPWR VPWR fd._2969_
+ sky130_fd_sc_hd__o31a_1
XFILLER_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7063_ fd._1304_ fd._2294_ VGND VGND VPWR VPWR fd._2296_ sky130_fd_sc_hd__nor2_1
Xfd._4275_ fd._2155_ fd._2188_ VGND VGND VPWR VPWR fd._2210_ sky130_fd_sc_hd__and2_1
XFILLER_81_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_82 VGND VGND VPWR VPWR user_project_wrapper_82/HI io_oeb[4]
+ sky130_fd_sc_hd__conb_1
Xuser_project_wrapper_93 VGND VGND VPWR VPWR user_project_wrapper_93/HI io_oeb[15]
+ sky130_fd_sc_hd__conb_1
XFILLER_228_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6014_ fd._0964_ VGND VGND VPWR VPWR fd._1142_ sky130_fd_sc_hd__inv_2
XFILLER_250_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7965_ fd._3174_ fd._3163_ fd._3173_ VGND VGND VPWR VPWR fd._3289_ sky130_fd_sc_hd__and3_1
XFILLER_52_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6916_ fd._0928_ VGND VGND VPWR VPWR fd._2135_ sky130_fd_sc_hd__buf_6
XFILLER_276_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7896_ fd._3081_ fd._3087_ fd._3212_ VGND VGND VPWR VPWR fd._3213_ sky130_fd_sc_hd__or3_1
XFILLER_50_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6847_ fd._1852_ fd._2058_ VGND VGND VPWR VPWR fd._2059_ sky130_fd_sc_hd__nand2_1
XFILLER_117_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6778_ fd._0450_ fd._1955_ VGND VGND VPWR VPWR fd._1983_ sky130_fd_sc_hd__nand2_1
XFILLER_137_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_1629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5729_ fd._0781_ fd._0794_ fd._0796_ fd._0800_ fd._3695_ VGND VGND VPWR VPWR fd._0829_
+ sky130_fd_sc_hd__a2111o_2
XFILLER_277_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_226_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_263_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_project_wrapper_109 VGND VGND VPWR VPWR user_project_wrapper_109/HI io_oeb[31]
+ sky130_fd_sc_hd__conb_1
XFILLER_110_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_272_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput43 net43 VGND VGND VPWR VPWR io_out[18] sky130_fd_sc_hd__buf_2
XTAP_6000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_218_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput54 net54 VGND VGND VPWR VPWR io_out[28] sky130_fd_sc_hd__buf_2
XTAP_6011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput65 net65 VGND VGND VPWR VPWR io_out[9] sky130_fd_sc_hd__buf_2
XFILLER_150_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_1584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_249_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_264_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_264_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_281_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7750_ fd._0768_ fd._3042_ fd._3048_ VGND VGND VPWR VPWR fd._3052_ sky130_fd_sc_hd__o21ai_1
XFILLER_9_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4962_ fd._4056_ fd._3919_ VGND VGND VPWR VPWR fd._4057_ sky130_fd_sc_hd__nand2_1
XFILLER_145_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6701_ fd._1856_ fd._1897_ VGND VGND VPWR VPWR fd._1898_ sky130_fd_sc_hd__xnor2_1
Xfd._7681_ fd._2965_ fd._2971_ fd._2972_ fd._2973_ fd._2975_ VGND VGND VPWR VPWR fd._2976_
+ sky130_fd_sc_hd__a2111o_1
Xfd._4893_ fd._3860_ fd._3986_ fd._3959_ VGND VGND VPWR VPWR fd._3987_ sky130_fd_sc_hd__mux2_1
XFILLER_184_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6632_ fd._1802_ fd._1804_ VGND VGND VPWR VPWR fd._1822_ sky130_fd_sc_hd__xnor2_1
XFILLER_12_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_259_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6563_ fd._1744_ fd._1745_ VGND VGND VPWR VPWR fd._1746_ sky130_fd_sc_hd__nand2_1
XFILLER_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5514_ fd._0585_ fd._0590_ fd._0591_ VGND VGND VPWR VPWR fd._0592_ sky130_fd_sc_hd__o21ai_2
XFILLER_141_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_1624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6494_ fd._1470_ fd._1669_ VGND VGND VPWR VPWR fd._1670_ sky130_fd_sc_hd__xnor2_1
XFILLER_140_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._8233_ net67 net18 VGND VGND VPWR VPWR fd.a\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_267_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5445_ fd._0507_ fd._0515_ VGND VGND VPWR VPWR fd._0517_ sky130_fd_sc_hd__nand2_1
XFILLER_79_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8164_ fd._3476_ fd._3477_ VGND VGND VPWR VPWR fd._3478_ sky130_fd_sc_hd__nand2_1
XFILLER_283_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5376_ fd._0258_ fd._0440_ VGND VGND VPWR VPWR fd._0441_ sky130_fd_sc_hd__or2_1
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7115_ fd._2157_ fd._2352_ fd._2322_ VGND VGND VPWR VPWR fd._2354_ sky130_fd_sc_hd__mux2_1
XFILLER_110_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4327_ fd._2749_ fd._2771_ VGND VGND VPWR VPWR fd._2782_ sky130_fd_sc_hd__xnor2_1
XFILLER_254_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8095_ fd._0651_ fd._0849_ fd._3411_ VGND VGND VPWR VPWR fd._3417_ sky130_fd_sc_hd__mux2_1
XFILLER_270_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7046_ fd._2270_ fd._2275_ fd._2277_ VGND VGND VPWR VPWR fd._2278_ sky130_fd_sc_hd__a21oi_1
XFILLER_74_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4258_ fd._1891_ fd._1935_ fd._2001_ fd._2012_ VGND VGND VPWR VPWR fd._2023_ sky130_fd_sc_hd__a31o_1
XFILLER_208_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4189_ fd._1253_ VGND VGND VPWR VPWR fd._1264_ sky130_fd_sc_hd__buf_6
XFILLER_223_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7948_ fd._2751_ fd._3267_ fd._3240_ fd._3269_ VGND VGND VPWR VPWR fd._3270_ sky130_fd_sc_hd__a211o_1
XFILLER_202_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_8908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7879_ fd._3191_ fd._3193_ fd._3076_ VGND VGND VPWR VPWR fd._3194_ sky130_fd_sc_hd__mux2_1
XFILLER_30_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_259_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_270_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5230_ fd._0271_ fd._0279_ VGND VGND VPWR VPWR fd._0280_ sky130_fd_sc_hd__nor2_1
XTAP_5173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_264_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5161_ fd._0201_ fd._0203_ VGND VGND VPWR VPWR fd._0204_ sky130_fd_sc_hd__xnor2_1
XTAP_4483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4112_ fd._0208_ fd._0285_ fd._0307_ fd._0406_ VGND VGND VPWR VPWR fd._0417_ sky130_fd_sc_hd__nand4bb_2
XFILLER_280_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5092_ fd._0050_ fd._0052_ fd._0057_ fd._0127_ VGND VGND VPWR VPWR fd._0128_ sky130_fd_sc_hd__a31o_1
XFILLER_45_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_251_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_260_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7802_ fd._2988_ fd._3107_ fd._3076_ fd._3108_ VGND VGND VPWR VPWR fd._3109_ sky130_fd_sc_hd__a31oi_1
XFILLER_192_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5994_ fd._0949_ fd._1119_ VGND VGND VPWR VPWR fd._1120_ sky130_fd_sc_hd__nand2_1
XFILLER_285_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7733_ fd._3027_ fd._3032_ fd._2877_ VGND VGND VPWR VPWR fd._3033_ sky130_fd_sc_hd__mux2_1
Xfd._4945_ fd._3716_ fd._4038_ VGND VGND VPWR VPWR fd._4039_ sky130_fd_sc_hd__or2_1
XFILLER_220_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7664_ fd._2763_ fd._2956_ VGND VGND VPWR VPWR fd._2957_ sky130_fd_sc_hd__and2_1
Xfd._4876_ fd._3969_ VGND VGND VPWR VPWR fd._3970_ sky130_fd_sc_hd__clkinv_2
XFILLER_172_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6615_ fd._1637_ fd._1710_ VGND VGND VPWR VPWR fd._1804_ sky130_fd_sc_hd__and2_1
XFILLER_86_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7595_ fd._2682_ fd._2820_ VGND VGND VPWR VPWR fd._2882_ sky130_fd_sc_hd__or2_1
XFILLER_141_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_259_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6546_ fd._1597_ fd._1727_ fd._1719_ VGND VGND VPWR VPWR fd._1728_ sky130_fd_sc_hd__mux2_1
XFILLER_87_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6477_ fd._1456_ fd._1651_ VGND VGND VPWR VPWR fd._1652_ sky130_fd_sc_hd__xnor2_1
XFILLER_101_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8216_ net72 net31 VGND VGND VPWR VPWR fd.a\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_228_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5428_ fd._0338_ fd._0336_ VGND VGND VPWR VPWR fd._0498_ sky130_fd_sc_hd__or2b_1
XFILLER_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_270_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8147_ fd._3460_ fd._3461_ VGND VGND VPWR VPWR fd._3462_ sky130_fd_sc_hd__nor2_1
Xfd._5359_ fd._0421_ fd._0235_ fd._0062_ VGND VGND VPWR VPWR fd._0422_ sky130_fd_sc_hd__mux2_1
XFILLER_215_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_270_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8078_ fd._2238_ fd._2423_ fd._3398_ VGND VGND VPWR VPWR fd._3406_ sky130_fd_sc_hd__mux2_1
XFILLER_262_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7029_ fd._2075_ fd._2102_ VGND VGND VPWR VPWR fd._2259_ sky130_fd_sc_hd__xor2_1
XFILLER_54_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_260_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_278_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_278_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_265_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_1576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_259_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_259_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4730_ fd._3732_ fd._3731_ VGND VGND VPWR VPWR fd._3824_ sky130_fd_sc_hd__and2b_1
XFILLER_185_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4661_ fd._3587_ fd._3754_ fd._3626_ VGND VGND VPWR VPWR fd._3755_ sky130_fd_sc_hd__mux2_1
XFILLER_29_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6400_ fd._1398_ fd._1400_ VGND VGND VPWR VPWR fd._1567_ sky130_fd_sc_hd__and2_1
XFILLER_83_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7380_ fd._2427_ fd._2644_ VGND VGND VPWR VPWR fd._2645_ sky130_fd_sc_hd__or2_1
XFILLER_116_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._4592_ fd._3534_ fd._3685_ fd._3624_ VGND VGND VPWR VPWR fd._3686_ sky130_fd_sc_hd__mux2_1
XFILLER_151_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6331_ fd._1490_ VGND VGND VPWR VPWR fd._1491_ sky130_fd_sc_hd__clkinv_4
XFILLER_116_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_270_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6262_ fd._0916_ fd._1350_ VGND VGND VPWR VPWR fd._1415_ sky130_fd_sc_hd__and2_1
XFILLER_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_285_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_1504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8001_ fd._3135_ fd._3314_ VGND VGND VPWR VPWR fd._3328_ sky130_fd_sc_hd__xnor2_1
XFILLER_49_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_266_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5213_ fd._3869_ fd._0240_ fd._0250_ VGND VGND VPWR VPWR fd._0261_ sky130_fd_sc_hd__and3_1
XFILLER_225_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6193_ fd._1338_ VGND VGND VPWR VPWR fd._1339_ sky130_fd_sc_hd__inv_2
XTAP_4280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_266_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5144_ fd._4059_ fd._0067_ VGND VGND VPWR VPWR fd._0185_ sky130_fd_sc_hd__nand2_1
XFILLER_64_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5075_ fd._4000_ fd._4004_ VGND VGND VPWR VPWR fd._0110_ sky130_fd_sc_hd__nand2_1
XFILLER_221_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_277_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5977_ fd._3905_ VGND VGND VPWR VPWR fd._1102_ sky130_fd_sc_hd__buf_6
XFILLER_277_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4928_ fd._4020_ fd._4021_ VGND VGND VPWR VPWR fd._4022_ sky130_fd_sc_hd__xor2_1
XFILLER_175_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7716_ fd._2055_ fd._3014_ VGND VGND VPWR VPWR fd._3015_ sky130_fd_sc_hd__nor2_1
XFILLER_12_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_259_1690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7647_ fd._2758_ fd._2767_ VGND VGND VPWR VPWR fd._2939_ sky130_fd_sc_hd__or2b_1
XFILLER_133_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4859_ fd._3946_ fd._3952_ VGND VGND VPWR VPWR fd._3953_ sky130_fd_sc_hd__or2b_1
XFILLER_47_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_270 VGND VGND VPWR VPWR user_project_wrapper_270/HI wbs_dat_o[16]
+ sky130_fd_sc_hd__conb_1
XFILLER_86_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_project_wrapper_281 VGND VGND VPWR VPWR user_project_wrapper_281/HI wbs_dat_o[27]
+ sky130_fd_sc_hd__conb_1
XFILLER_251_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7578_ fd._1816_ VGND VGND VPWR VPWR fd._2863_ sky130_fd_sc_hd__buf_6
XFILLER_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6529_ fd._1304_ fd._1708_ VGND VGND VPWR VPWR fd._1709_ sky130_fd_sc_hd__nor2_1
XFILLER_141_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_284_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_279_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5900_ fd._1016_ fd._0831_ VGND VGND VPWR VPWR fd._1017_ sky130_fd_sc_hd__and2b_1
XFILLER_141_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._6880_ fd._2084_ fd._2088_ fd._2092_ fd._2094_ VGND VGND VPWR VPWR fd._2095_ sky130_fd_sc_hd__o211a_1
XFILLER_159_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5831_ fd._3905_ fd._0938_ VGND VGND VPWR VPWR fd._0941_ sky130_fd_sc_hd__and2_1
XFILLER_200_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_278_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5762_ fd._0779_ fd._0763_ VGND VGND VPWR VPWR fd._0865_ sky130_fd_sc_hd__or2b_1
XFILLER_183_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7501_ fd._2777_ VGND VGND VPWR VPWR fd._2778_ sky130_fd_sc_hd__clkinv_4
Xfd._4713_ fd._3806_ fd._3636_ fd._3788_ VGND VGND VPWR VPWR fd._3807_ sky130_fd_sc_hd__mux2_1
XFILLER_170_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5693_ fd._0786_ fd._0788_ VGND VGND VPWR VPWR fd._0789_ sky130_fd_sc_hd__nand2_1
XFILLER_131_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7432_ fd._2700_ fd._2677_ fd._2701_ VGND VGND VPWR VPWR fd._2702_ sky130_fd_sc_hd__a21oi_2
Xfd._4644_ fd._3646_ fd._3733_ fd._3737_ VGND VGND VPWR VPWR fd._3738_ sky130_fd_sc_hd__mux2_1
XFILLER_215_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_272_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7363_ fd._2623_ fd._2625_ VGND VGND VPWR VPWR fd._2626_ sky130_fd_sc_hd__nand2_1
XFILLER_123_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4575_ fd.b\[6\] VGND VGND VPWR VPWR fd._3669_ sky130_fd_sc_hd__buf_6
XFILLER_215_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_250_1440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_284_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6314_ fd._1471_ VGND VGND VPWR VPWR fd._1472_ sky130_fd_sc_hd__clkinv_2
XFILLER_22_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7294_ fd._2546_ fd._2549_ fd._2505_ VGND VGND VPWR VPWR fd._2550_ sky130_fd_sc_hd__mux2_1
XFILLER_244_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6245_ fd._0638_ VGND VGND VPWR VPWR fd._1397_ sky130_fd_sc_hd__buf_6
XFILLER_49_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_285_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6176_ fd._1317_ fd._1320_ fd._1232_ VGND VGND VPWR VPWR fd._1321_ sky130_fd_sc_hd__mux2_1
XFILLER_65_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5127_ fd._0079_ fd._0165_ VGND VGND VPWR VPWR fd._0167_ sky130_fd_sc_hd__nor2_1
XFILLER_94_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5058_ fd._0083_ fd._0088_ fd._0090_ VGND VGND VPWR VPWR fd._0091_ sky130_fd_sc_hd__a21o_1
XFILLER_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_256_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_256_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_263_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_1686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_9044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_9055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_285_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4360_ fd._2738_ fd._2793_ VGND VGND VPWR VPWR fd._3145_ sky130_fd_sc_hd__nand2_1
XTAP_6996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_281_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4291_ fd.b\[13\] fd._1429_ VGND VGND VPWR VPWR fd._2386_ sky130_fd_sc_hd__and2_1
XFILLER_130_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6030_ fd._0207_ fd._1159_ VGND VGND VPWR VPWR fd._1160_ sky130_fd_sc_hd__xnor2_1
XFILLER_62_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._7981_ fd._1751_ fd._3286_ fd._3291_ fd._2533_ VGND VGND VPWR VPWR fd._3306_ sky130_fd_sc_hd__o22a_1
XFILLER_280_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6932_ fd._2150_ fd._2151_ VGND VGND VPWR VPWR fd._2152_ sky130_fd_sc_hd__or2_1
XFILLER_147_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6863_ fd._0726_ VGND VGND VPWR VPWR fd._2076_ sky130_fd_sc_hd__buf_6
XFILLER_147_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5814_ fd._0680_ fd._0921_ fd._0801_ VGND VGND VPWR VPWR fd._0922_ sky130_fd_sc_hd__mux2_1
XFILLER_200_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6794_ fd._1998_ fd._1999_ fd._1969_ VGND VGND VPWR VPWR fd._2000_ sky130_fd_sc_hd__a21oi_1
XFILLER_116_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5745_ fd._0845_ VGND VGND VPWR VPWR fd._0847_ sky130_fd_sc_hd__clkinv_2
XFILLER_176_1647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_1379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5676_ fd._0767_ fd._0770_ VGND VGND VPWR VPWR fd._0771_ sky130_fd_sc_hd__and2_1
XFILLER_276_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_252_1546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4627_ fd._3716_ fd._3720_ VGND VGND VPWR VPWR fd._3721_ sky130_fd_sc_hd__nor2_1
XFILLER_252_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7415_ fd._2682_ VGND VGND VPWR VPWR fd._2684_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_217_1688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7346_ fd._2601_ fd._2605_ fd._2607_ VGND VGND VPWR VPWR fd._2608_ sky130_fd_sc_hd__o21ai_1
XFILLER_135_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4558_ fd._3548_ fd._3647_ VGND VGND VPWR VPWR fd._3652_ sky130_fd_sc_hd__xnor2_1
XFILLER_97_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_242_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7277_ fd._2531_ VGND VGND VPWR VPWR fd._2532_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_284_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4489_ fd._3582_ VGND VGND VPWR VPWR fd._3583_ sky130_fd_sc_hd__clkinv_4
XFILLER_66_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6228_ fd._0821_ fd._1210_ fd._1212_ VGND VGND VPWR VPWR fd._1378_ sky130_fd_sc_hd__a21o_1
XFILLER_81_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_253_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6159_ fd._0207_ fd._1301_ VGND VGND VPWR VPWR fd._1302_ sky130_fd_sc_hd__xnor2_1
XFILLER_164_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_1670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_283_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_251_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_270_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_268_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_262_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_275_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_279_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_7 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5530_ fd._0480_ fd._0609_ VGND VGND VPWR VPWR fd._0610_ sky130_fd_sc_hd__nand2_1
XFILLER_193_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_273_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5461_ fd._0533_ VGND VGND VPWR VPWR fd._0534_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_136_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7200_ fd._2446_ VGND VGND VPWR VPWR fd._2447_ sky130_fd_sc_hd__inv_2
XFILLER_117_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4412_ fd._3503_ fd._3505_ VGND VGND VPWR VPWR fd._3506_ sky130_fd_sc_hd__xnor2_1
XTAP_6771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8180_ net77 fd.mc\[4\] VGND VGND VPWR VPWR fd.c\[4\] sky130_fd_sc_hd__dfxtp_1
Xfd._5392_ fd._0419_ fd._0457_ VGND VGND VPWR VPWR fd._0458_ sky130_fd_sc_hd__xnor2_1
XTAP_6793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7131_ fd._2184_ fd._2370_ VGND VGND VPWR VPWR fd._2371_ sky130_fd_sc_hd__and2_1
Xfd._4343_ fd.b\[19\] fd._2914_ VGND VGND VPWR VPWR fd._2958_ sky130_fd_sc_hd__or2_1
XFILLER_266_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7062_ fd._1304_ fd._2294_ VGND VGND VPWR VPWR fd._2295_ sky130_fd_sc_hd__nand2_1
XFILLER_63_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4274_ fd._2155_ fd._2188_ VGND VGND VPWR VPWR fd._2199_ sky130_fd_sc_hd__nor2_1
XFILLER_130_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6013_ fd._0963_ VGND VGND VPWR VPWR fd._1141_ sky130_fd_sc_hd__clkinv_2
XFILLER_282_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_83 VGND VGND VPWR VPWR user_project_wrapper_83/HI io_oeb[5]
+ sky130_fd_sc_hd__conb_1
Xuser_project_wrapper_94 VGND VGND VPWR VPWR user_project_wrapper_94/HI io_oeb[16]
+ sky130_fd_sc_hd__conb_1
XFILLER_179_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_250_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_280_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7964_ fd._3158_ VGND VGND VPWR VPWR fd._3287_ sky130_fd_sc_hd__clkinv_2
XFILLER_241_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6915_ fd._2131_ fd._2132_ VGND VGND VPWR VPWR fd._2134_ sky130_fd_sc_hd__or2_1
XFILLER_223_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._7895_ fd._3093_ fd._3096_ fd._3207_ fd._3208_ fd._3210_ VGND VGND VPWR VPWR fd._3212_
+ sky130_fd_sc_hd__a311oi_1
XFILLER_50_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6846_ fd._1494_ fd._1851_ VGND VGND VPWR VPWR fd._2058_ sky130_fd_sc_hd__or2_1
XFILLER_239_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6777_ fd._1958_ fd._1965_ fd._1975_ fd._1981_ VGND VGND VPWR VPWR fd._1982_ sky130_fd_sc_hd__o211a_1
XFILLER_117_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5728_ fd._0820_ fd._0827_ VGND VGND VPWR VPWR fd._0828_ sky130_fd_sc_hd__and2_1
XFILLER_277_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5659_ fd._0585_ fd._0751_ VGND VGND VPWR VPWR fd._0752_ sky130_fd_sc_hd__xnor2_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7329_ fd._2335_ fd._2588_ VGND VGND VPWR VPWR fd._2589_ sky130_fd_sc_hd__xnor2_1
XTAP_3419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_1685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_272_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_263_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_263_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput44 net44 VGND VGND VPWR VPWR io_out[19] sky130_fd_sc_hd__buf_2
XTAP_6001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput55 net55 VGND VGND VPWR VPWR io_out[29] sky130_fd_sc_hd__buf_2
XTAP_6023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_264_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_1670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_281_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_1523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_1518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._4961_ fd._3841_ fd._3916_ fd._3839_ VGND VGND VPWR VPWR fd._4056_ sky130_fd_sc_hd__a21o_1
XFILLER_185_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6700_ fd._1864_ fd._1892_ fd._1895_ fd._1896_ VGND VGND VPWR VPWR fd._1897_ sky130_fd_sc_hd__o31a_1
XFILLER_8_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7680_ fd._2918_ fd._2974_ VGND VGND VPWR VPWR fd._2975_ sky130_fd_sc_hd__nand2_1
Xfd._4892_ fd._3984_ fd._3985_ VGND VGND VPWR VPWR fd._3986_ sky130_fd_sc_hd__xor2_1
XFILLER_199_1499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_275_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6631_ fd._1810_ fd._1811_ fd._1815_ fd._1820_ VGND VGND VPWR VPWR fd._1821_ sky130_fd_sc_hd__a22oi_4
XFILLER_201_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6562_ fd._1178_ fd._1743_ VGND VGND VPWR VPWR fd._1745_ sky130_fd_sc_hd__or2_1
XFILLER_154_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5513_ fd._1264_ fd._0589_ VGND VGND VPWR VPWR fd._0591_ sky130_fd_sc_hd__nand2_1
XFILLER_140_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6493_ fd._1476_ fd._1475_ VGND VGND VPWR VPWR fd._1669_ sky130_fd_sc_hd__nor2_1
XFILLER_86_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_1674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8232_ net66 net17 VGND VGND VPWR VPWR fd.a\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_234_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5444_ fd._0324_ fd._0325_ VGND VGND VPWR VPWR fd._0515_ sky130_fd_sc_hd__nand2_1
XFILLER_214_1647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_214_1669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8163_ fd.a\[29\] fd.b\[29\] VGND VGND VPWR VPWR fd._3477_ sky130_fd_sc_hd__or2b_1
XFILLER_227_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5375_ fd._4011_ fd._3689_ fd._0242_ fd._0244_ VGND VGND VPWR VPWR fd._0440_ sky130_fd_sc_hd__and4_1
XFILLER_223_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._7114_ fd._2350_ fd._2351_ VGND VGND VPWR VPWR fd._2352_ sky130_fd_sc_hd__xnor2_1
XFILLER_269_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4326_ fd._2760_ fd._1154_ VGND VGND VPWR VPWR fd._2771_ sky130_fd_sc_hd__nor2_1
XFILLER_48_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8094_ fd._3415_ VGND VGND VPWR VPWR fd.mc\[14\] sky130_fd_sc_hd__clkbuf_1
XFILLER_247_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_242_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7045_ fd._0382_ fd._2274_ VGND VGND VPWR VPWR fd._2277_ sky130_fd_sc_hd__nor2_1
Xfd._4257_ fd.b\[3\] fd._1880_ VGND VGND VPWR VPWR fd._2012_ sky130_fd_sc_hd__nor2_1
XFILLER_169_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_251_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4188_ fd.b\[17\] VGND VGND VPWR VPWR fd._1253_ sky130_fd_sc_hd__buf_6
XFILLER_211_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7947_ fd._3268_ VGND VGND VPWR VPWR fd._3269_ sky130_fd_sc_hd__inv_2
XFILLER_109_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_276_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7878_ fd._3192_ fd._2972_ VGND VGND VPWR VPWR fd._3193_ sky130_fd_sc_hd__xnor2_1
XFILLER_258_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6829_ fd._1842_ fd._1907_ VGND VGND VPWR VPWR fd._2039_ sky130_fd_sc_hd__or2_1
XFILLER_85_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_254_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_277_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_264_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_218_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_249_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5160_ fd._0202_ fd._0007_ VGND VGND VPWR VPWR fd._0203_ sky130_fd_sc_hd__nor2_1
XTAP_4473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4111_ fd._0318_ fd.a\[3\] fd._0351_ fd._0395_ fd._0329_ VGND VGND VPWR VPWR fd._0406_
+ sky130_fd_sc_hd__a221o_1
XFILLER_218_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5091_ fd._4011_ fd._0122_ VGND VGND VPWR VPWR fd._0127_ sky130_fd_sc_hd__xnor2_1
XTAP_3783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7801_ fd._2898_ fd._3076_ VGND VGND VPWR VPWR fd._3108_ sky130_fd_sc_hd__nor2_1
XFILLER_140_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5993_ fd._0942_ fd._0947_ fd._0951_ VGND VGND VPWR VPWR fd._1119_ sky130_fd_sc_hd__a21o_1
XFILLER_185_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._7732_ fd._3031_ fd._2846_ VGND VGND VPWR VPWR fd._3032_ sky130_fd_sc_hd__xor2_1
XFILLER_9_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4944_ fd._3903_ fd._4037_ fd._3960_ VGND VGND VPWR VPWR fd._4038_ sky130_fd_sc_hd__mux2_1
XFILLER_51_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4875_ fd._3968_ fd._3925_ VGND VGND VPWR VPWR fd._3969_ sky130_fd_sc_hd__xor2_1
Xfd._7663_ fd._2953_ fd._2955_ fd._2874_ VGND VGND VPWR VPWR fd._2956_ sky130_fd_sc_hd__mux2_1
XFILLER_12_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6614_ fd._1703_ fd._1709_ fd._1717_ VGND VGND VPWR VPWR fd._1802_ sky130_fd_sc_hd__o21ai_1
XFILLER_216_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._7594_ fd._2679_ VGND VGND VPWR VPWR fd._2880_ sky130_fd_sc_hd__clkinv_2
XFILLER_86_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_259_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6545_ fd._1723_ fd._1725_ VGND VGND VPWR VPWR fd._1727_ sky130_fd_sc_hd__xnor2_1
XFILLER_173_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._6476_ fd._1457_ fd._1458_ VGND VGND VPWR VPWR fd._1651_ sky130_fd_sc_hd__nand2_1
XFILLER_228_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_268_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_267_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8215_ net72 net30 VGND VGND VPWR VPWR fd.a\[7\] sky130_fd_sc_hd__dfxtp_1
Xfd._5427_ fd._0335_ VGND VGND VPWR VPWR fd._0497_ sky130_fd_sc_hd__clkinv_2
XFILLER_110_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_283_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_283_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5358_ fd._0239_ fd._0235_ VGND VGND VPWR VPWR fd._0421_ sky130_fd_sc_hd__nand2_1
Xfd._8146_ fd.a\[27\] fd.b\[27\] VGND VGND VPWR VPWR fd._3461_ sky130_fd_sc_hd__and2b_1
XFILLER_103_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4309_ fd.b\[16\] VGND VGND VPWR VPWR fd._2584_ sky130_fd_sc_hd__buf_6
XFILLER_110_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8077_ fd._3405_ VGND VGND VPWR VPWR fd.mc\[6\] sky130_fd_sc_hd__clkbuf_1
Xfd._5289_ fd._0146_ fd._0293_ fd._0088_ VGND VGND VPWR VPWR fd._0345_ sky130_fd_sc_hd__o21a_1
XFILLER_184_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7028_ fd._2256_ fd._2257_ VGND VGND VPWR VPWR fd._2258_ sky130_fd_sc_hd__nor2_1
XFILLER_251_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_1540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_221_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_275_74 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_1588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_267_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_259_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4660_ fd._3753_ fd._3593_ VGND VGND VPWR VPWR fd._3754_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4591_ fd._3538_ fd._3684_ VGND VGND VPWR VPWR fd._3685_ sky130_fd_sc_hd__xnor2_1
XFILLER_190_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6330_ fd._1444_ fd._1489_ VGND VGND VPWR VPWR fd._1490_ sky130_fd_sc_hd__and2_1
XFILLER_155_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6261_ fd._1361_ fd._1413_ fd._1359_ VGND VGND VPWR VPWR fd._1414_ sky130_fd_sc_hd__a21oi_1
XFILLER_265_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5212_ fd._0257_ fd._0259_ VGND VGND VPWR VPWR fd._0260_ sky130_fd_sc_hd__nor2_1
Xfd._8000_ fd._1173_ fd._3326_ VGND VGND VPWR VPWR fd._3327_ sky130_fd_sc_hd__nor2_1
XFILLER_264_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_265_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6192_ fd._1304_ fd._1306_ VGND VGND VPWR VPWR fd._1338_ sky130_fd_sc_hd__and2_1
XFILLER_266_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5143_ fd._4054_ fd._4061_ VGND VGND VPWR VPWR fd._0184_ sky130_fd_sc_hd__nor2_1
XFILLER_280_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5074_ fd._0106_ fd._0107_ VGND VGND VPWR VPWR fd._0108_ sky130_fd_sc_hd__xnor2_1
XFILLER_233_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5976_ fd._3905_ fd._1100_ VGND VGND VPWR VPWR fd._1101_ sky130_fd_sc_hd__nor2_1
XFILLER_146_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_277_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7715_ fd._3012_ VGND VGND VPWR VPWR fd._3014_ sky130_fd_sc_hd__clkinvlp_2
Xfd._4927_ fd._3862_ fd._3885_ VGND VGND VPWR VPWR fd._4021_ sky130_fd_sc_hd__and2_1
XFILLER_161_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_255_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7646_ fd._2764_ fd._2766_ VGND VGND VPWR VPWR fd._2938_ sky130_fd_sc_hd__or2_1
Xfd._4858_ fd._3950_ fd._3951_ VGND VGND VPWR VPWR fd._3952_ sky130_fd_sc_hd__nor2_1
XFILLER_245_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_project_wrapper_260 VGND VGND VPWR VPWR user_project_wrapper_260/HI wbs_dat_o[6]
+ sky130_fd_sc_hd__conb_1
XFILLER_47_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_271 VGND VGND VPWR VPWR user_project_wrapper_271/HI wbs_dat_o[17]
+ sky130_fd_sc_hd__conb_1
XFILLER_88_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_282 VGND VGND VPWR VPWR user_project_wrapper_282/HI wbs_dat_o[28]
+ sky130_fd_sc_hd__conb_1
XFILLER_86_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7577_ fd._1816_ fd._2861_ VGND VGND VPWR VPWR fd._2862_ sky130_fd_sc_hd__and2_1
Xfd._4789_ fd._0252_ VGND VGND VPWR VPWR fd._3883_ sky130_fd_sc_hd__buf_6
XFILLER_141_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6528_ fd._1433_ fd._1707_ fd._1617_ VGND VGND VPWR VPWR fd._1708_ sky130_fd_sc_hd__mux2_1
XFILLER_29_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6459_ fd._1088_ VGND VGND VPWR VPWR fd._1632_ sky130_fd_sc_hd__buf_2
XFILLER_25_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_255_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_270_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8129_ fd._3442_ fd._3443_ VGND VGND VPWR VPWR fd._3444_ sky130_fd_sc_hd__nor2_1
XFILLER_215_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_1657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_260_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_279_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_279_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5830_ fd._0939_ VGND VGND VPWR VPWR fd._0940_ sky130_fd_sc_hd__inv_2
XFILLER_278_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5761_ fd._0755_ fd._0756_ VGND VGND VPWR VPWR fd._0864_ sky130_fd_sc_hd__nand2_1
XFILLER_170_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7500_ fd._2135_ fd._2776_ VGND VGND VPWR VPWR fd._2777_ sky130_fd_sc_hd__nand2_1
XFILLER_13_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4712_ fd._3804_ fd._3805_ VGND VGND VPWR VPWR fd._3806_ sky130_fd_sc_hd__or2_1
Xfd._5692_ fd._0468_ fd._0787_ fd._0651_ VGND VGND VPWR VPWR fd._0788_ sky130_fd_sc_hd__mux2_1
XFILLER_87_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7431_ fd._2598_ fd._2670_ fd._2675_ VGND VGND VPWR VPWR fd._2701_ sky130_fd_sc_hd__and3_1
Xfd._4643_ fd._3734_ fd._3736_ VGND VGND VPWR VPWR fd._3737_ sky130_fd_sc_hd__xnor2_1
XFILLER_130_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_285_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._4574_ fd.b\[6\] fd._3667_ VGND VGND VPWR VPWR fd._3668_ sky130_fd_sc_hd__or2_1
Xfd._7362_ fd._2624_ fd._2489_ VGND VGND VPWR VPWR fd._2625_ sky130_fd_sc_hd__xnor2_1
XFILLER_96_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6313_ fd._1248_ fd._1276_ VGND VGND VPWR VPWR fd._1471_ sky130_fd_sc_hd__xnor2_1
XFILLER_250_1463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7293_ fd._2381_ fd._2548_ VGND VGND VPWR VPWR fd._2549_ sky130_fd_sc_hd__xnor2_1
XFILLER_250_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6244_ fd._1340_ fd._1348_ fd._1394_ fd._1384_ VGND VGND VPWR VPWR fd._1395_ sky130_fd_sc_hd__a22oi_2
XFILLER_285_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_237_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_252_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6175_ fd._1318_ fd._1071_ VGND VGND VPWR VPWR fd._1320_ sky130_fd_sc_hd__xnor2_1
XFILLER_64_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5126_ fd._0079_ fd._0165_ VGND VGND VPWR VPWR fd._0166_ sky130_fd_sc_hd__xor2_1
XFILLER_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5057_ fd._0089_ fd._0082_ VGND VGND VPWR VPWR fd._0090_ sky130_fd_sc_hd__and2_1
XFILLER_221_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5959_ fd._0908_ fd._1081_ fd._1046_ VGND VGND VPWR VPWR fd._1082_ sky130_fd_sc_hd__mux2_1
XFILLER_146_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_277_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7629_ fd._2566_ fd._2911_ VGND VGND VPWR VPWR fd._2919_ sky130_fd_sc_hd__and2_1
XFILLER_47_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_276_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_275_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_276_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_271_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_262_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_262_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_281_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4290_ fd._1627_ fd._2320_ fd._2353_ fd._2364_ VGND VGND VPWR VPWR fd._2375_ sky130_fd_sc_hd__a211o_1
XFILLER_219_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_281_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_267_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7980_ fd._3298_ fd._3303_ fd._3304_ VGND VGND VPWR VPWR fd._3305_ sky130_fd_sc_hd__or3b_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6931_ fd._2141_ fd._2149_ VGND VGND VPWR VPWR fd._2151_ sky130_fd_sc_hd__nor2_1
XFILLER_163_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6862_ fd._2073_ fd._2074_ VGND VGND VPWR VPWR fd._2075_ sky130_fd_sc_hd__nand2_1
XFILLER_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5813_ fd._0682_ fd._0920_ VGND VGND VPWR VPWR fd._0921_ sky130_fd_sc_hd__xnor2_1
XFILLER_162_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6793_ fd._1729_ fd._1920_ fd._1785_ VGND VGND VPWR VPWR fd._1999_ sky130_fd_sc_hd__or3_1
XFILLER_155_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5744_ fd._0840_ fd._0792_ VGND VGND VPWR VPWR fd._0845_ sky130_fd_sc_hd__xnor2_1
XFILLER_115_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_256_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5675_ fd._0768_ fd._0766_ VGND VGND VPWR VPWR fd._0770_ sky130_fd_sc_hd__nand2_1
XFILLER_135_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_252_1536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7414_ fd._2680_ fd._2681_ VGND VGND VPWR VPWR fd._2682_ sky130_fd_sc_hd__and2_1
XFILLER_44_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4626_ fd._3552_ fd._3719_ VGND VGND VPWR VPWR fd._3720_ sky130_fd_sc_hd__xnor2_1
XFILLER_258_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_1678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_284_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7345_ fd._1666_ fd._2604_ VGND VGND VPWR VPWR fd._2607_ sky130_fd_sc_hd__or2_1
XFILLER_85_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4557_ fd._0857_ fd._3650_ VGND VGND VPWR VPWR fd._3651_ sky130_fd_sc_hd__nor2_1
XFILLER_57_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4488_ fd._3579_ fd._3581_ VGND VGND VPWR VPWR fd._3582_ sky130_fd_sc_hd__nand2_1
Xfd._7276_ fd._2141_ fd._2530_ VGND VGND VPWR VPWR fd._2531_ sky130_fd_sc_hd__xnor2_1
XFILLER_2_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_285_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6227_ fd._0807_ fd._1376_ VGND VGND VPWR VPWR fd._1377_ sky130_fd_sc_hd__nand2_1
XFILLER_148_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6158_ fd._1152_ fd._1300_ fd._1232_ VGND VGND VPWR VPWR fd._1301_ sky130_fd_sc_hd__mux2_1
XFILLER_81_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_263_1643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5109_ fd._0146_ VGND VGND VPWR VPWR fd._0147_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_146_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6089_ fd._1219_ fd._1224_ VGND VGND VPWR VPWR fd._1225_ sky130_fd_sc_hd__nor2_1
XFILLER_222_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_263_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_263_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_1503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_8 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_8130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_8196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5460_ fd._0526_ fd._0530_ VGND VGND VPWR VPWR fd._0533_ sky130_fd_sc_hd__nand2_1
XFILLER_45_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4411_ fd._1759_ fd._3504_ VGND VGND VPWR VPWR fd._3505_ sky130_fd_sc_hd__nand2_1
XTAP_6772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5391_ fd._0456_ fd._0411_ fd._0409_ VGND VGND VPWR VPWR fd._0457_ sky130_fd_sc_hd__o21ai_1
XFILLER_136_1698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_282_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4342_ fd._0021_ fd._2936_ fd._1220_ VGND VGND VPWR VPWR fd._2947_ sky130_fd_sc_hd__mux2_1
XFILLER_255_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7130_ fd._1976_ fd._2368_ VGND VGND VPWR VPWR fd._2370_ sky130_fd_sc_hd__nand2_1
XFILLER_212_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_282_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4273_ fd._0439_ fd._2177_ fd._1220_ VGND VGND VPWR VPWR fd._2188_ sky130_fd_sc_hd__mux2_1
XFILLER_235_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7061_ fd._2061_ fd._2293_ fd._2238_ VGND VGND VPWR VPWR fd._2294_ sky130_fd_sc_hd__mux2_1
XFILLER_47_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6012_ fd._1133_ fd._1138_ fd._1139_ VGND VGND VPWR VPWR fd._1140_ sky130_fd_sc_hd__a21o_1
XFILLER_21_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_84 VGND VGND VPWR VPWR user_project_wrapper_84/HI io_oeb[6]
+ sky130_fd_sc_hd__conb_1
XFILLER_228_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_95 VGND VGND VPWR VPWR user_project_wrapper_95/HI io_oeb[17]
+ sky130_fd_sc_hd__conb_1
XFILLER_250_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_280_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7963_ fd._3162_ fd._3285_ fd._3240_ VGND VGND VPWR VPWR fd._3286_ sky130_fd_sc_hd__mux2_1
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6914_ fd._1173_ fd._2129_ VGND VGND VPWR VPWR fd._2132_ sky130_fd_sc_hd__nor2_1
Xfd._7894_ fd._3087_ fd._3209_ VGND VGND VPWR VPWR fd._3210_ sky130_fd_sc_hd__or2_1
XFILLER_223_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6845_ fd._2055_ fd._1898_ fd._1899_ VGND VGND VPWR VPWR fd._2057_ sky130_fd_sc_hd__a21o_1
XFILLER_163_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6776_ fd._1976_ fd._1978_ fd._1980_ fd._1585_ VGND VGND VPWR VPWR fd._1981_ sky130_fd_sc_hd__a211o_1
XFILLER_116_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5727_ fd._0632_ fd._0631_ VGND VGND VPWR VPWR fd._0827_ sky130_fd_sc_hd__nand2_1
XFILLER_171_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_256_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5658_ fd._0750_ fd._0590_ VGND VGND VPWR VPWR fd._0751_ sky130_fd_sc_hd__nor2_1
XFILLER_115_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4609_ fd._3510_ fd._3656_ VGND VGND VPWR VPWR fd._3703_ sky130_fd_sc_hd__xnor2_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5589_ fd._0511_ fd._0614_ fd._0674_ VGND VGND VPWR VPWR fd._0675_ sky130_fd_sc_hd__o21a_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7328_ fd._2347_ fd._2398_ VGND VGND VPWR VPWR fd._2588_ sky130_fd_sc_hd__nor2_1
XFILLER_6_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7259_ fd._2389_ fd._2511_ VGND VGND VPWR VPWR fd._2512_ sky130_fd_sc_hd__xnor2_1
XFILLER_26_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_278_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_259_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_272_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput34 net34 VGND VGND VPWR VPWR io_out[0] sky130_fd_sc_hd__buf_2
XFILLER_268_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput45 net45 VGND VGND VPWR VPWR io_out[1] sky130_fd_sc_hd__buf_2
XFILLER_27_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput56 net56 VGND VGND VPWR VPWR io_out[2] sky130_fd_sc_hd__buf_2
XTAP_6024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_1499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_264_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._4960_ fd._3734_ VGND VGND VPWR VPWR fd._4055_ sky130_fd_sc_hd__buf_8
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._4891_ fd._3861_ fd._3884_ VGND VGND VPWR VPWR fd._3985_ sky130_fd_sc_hd__nor2_1
XFILLER_8_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6630_ fd._1816_ fd._1819_ VGND VGND VPWR VPWR fd._1820_ sky130_fd_sc_hd__nor2_1
XFILLER_201_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6561_ fd._1178_ fd._1743_ VGND VGND VPWR VPWR fd._1744_ sky130_fd_sc_hd__nand2_1
XFILLER_153_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_1629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5512_ fd._1264_ fd._0589_ VGND VGND VPWR VPWR fd._0590_ sky130_fd_sc_hd__nor2_1
XFILLER_158_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._6492_ fd._1659_ fd._1662_ fd._1665_ fd._1667_ VGND VGND VPWR VPWR fd._1668_ sky130_fd_sc_hd__a31oi_2
XFILLER_140_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8231_ net66 net16 VGND VGND VPWR VPWR fd.a\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_7292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5443_ fd._0512_ fd._0513_ VGND VGND VPWR VPWR fd._0514_ sky130_fd_sc_hd__nor2_1
XFILLER_79_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8162_ fd.b\[29\] fd.a\[29\] VGND VGND VPWR VPWR fd._3476_ sky130_fd_sc_hd__or2b_1
XFILLER_283_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5374_ fd._0437_ fd._0270_ VGND VGND VPWR VPWR fd._0438_ sky130_fd_sc_hd__nand2_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7113_ fd._2158_ fd._2191_ VGND VGND VPWR VPWR fd._2351_ sky130_fd_sc_hd__and2b_1
XFILLER_283_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4325_ fd._1165_ fd.a\[21\] VGND VGND VPWR VPWR fd._2760_ sky130_fd_sc_hd__nor2_1
XFILLER_236_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8093_ fd._0849_ fd._1047_ fd._3411_ VGND VGND VPWR VPWR fd._3415_ sky130_fd_sc_hd__mux2_1
XFILLER_130_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7044_ fd._0382_ fd._2274_ VGND VGND VPWR VPWR fd._2275_ sky130_fd_sc_hd__nand2_1
XFILLER_247_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._4256_ fd.b\[0\] fd._1968_ fd._1979_ fd._1990_ VGND VGND VPWR VPWR fd._2001_ sky130_fd_sc_hd__o211ai_1
XFILLER_165_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_235_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_251_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4187_ fd._1165_ VGND VGND VPWR VPWR fd._1242_ sky130_fd_sc_hd__buf_6
XFILLER_50_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_280_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7946_ fd._3077_ fd._3165_ fd._3168_ VGND VGND VPWR VPWR fd._3268_ sky130_fd_sc_hd__a21oi_1
XFILLER_17_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7877_ fd._2974_ fd._3181_ fd._2918_ VGND VGND VPWR VPWR fd._3192_ sky130_fd_sc_hd__a21bo_1
XFILLER_164_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6828_ fd._1848_ fd._1905_ VGND VGND VPWR VPWR fd._2038_ sky130_fd_sc_hd__nand2_1
XFILLER_117_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6759_ fd._1767_ fd._1960_ fd._1961_ VGND VGND VPWR VPWR fd._1962_ sky130_fd_sc_hd__and3_1
XFILLER_277_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_264_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_277_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_280_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1579 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_249_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_265_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_264_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4110_ fd._0362_ fd._0373_ fd._0384_ VGND VGND VPWR VPWR fd._0395_ sky130_fd_sc_hd__a21o_1
XFILLER_229_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5090_ fd._0059_ fd._0121_ fd._0124_ fd._0125_ VGND VGND VPWR VPWR fd._0126_ sky130_fd_sc_hd__a211o_1
XFILLER_166_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7800_ fd._2986_ fd._3106_ VGND VGND VPWR VPWR fd._3107_ sky130_fd_sc_hd__nand2_1
XFILLER_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5992_ fd._3917_ VGND VGND VPWR VPWR fd._1118_ sky130_fd_sc_hd__buf_6
XFILLER_146_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7731_ fd._3029_ fd._3030_ fd._2836_ VGND VGND VPWR VPWR fd._3031_ sky130_fd_sc_hd__o21a_1
XFILLER_8_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4943_ fd._4036_ fd._3907_ VGND VGND VPWR VPWR fd._4037_ sky130_fd_sc_hd__xnor2_1
XFILLER_146_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7662_ fd._2946_ fd._2954_ VGND VGND VPWR VPWR fd._2955_ sky130_fd_sc_hd__or2b_1
XFILLER_255_1704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._4874_ fd._3821_ fd._3923_ VGND VGND VPWR VPWR fd._3968_ sky130_fd_sc_hd__nand2_1
XFILLER_177_1551 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6613_ fd._1796_ fd._1800_ VGND VGND VPWR VPWR fd._1801_ sky130_fd_sc_hd__xnor2_1
XFILLER_114_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7593_ fd._2819_ fd._2822_ fd._2876_ fd._2878_ VGND VGND VPWR VPWR fd._2879_ sky130_fd_sc_hd__o31a_1
XFILLER_82_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_259_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6544_ fd._1724_ fd._1598_ VGND VGND VPWR VPWR fd._1725_ sky130_fd_sc_hd__nor2_1
XFILLER_253_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_259_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_275_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6475_ fd._1608_ fd._1610_ fd._1609_ VGND VGND VPWR VPWR fd._1650_ sky130_fd_sc_hd__o21bai_1
XFILLER_256_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8214_ net72 net29 VGND VGND VPWR VPWR fd.a\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_228_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5426_ fd._0089_ fd._0495_ VGND VGND VPWR VPWR fd._0496_ sky130_fd_sc_hd__or2_1
XFILLER_214_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8145_ fd.b\[27\] fd.a\[27\] VGND VGND VPWR VPWR fd._3460_ sky130_fd_sc_hd__and2b_1
Xfd._5357_ fd._0409_ fd._0418_ VGND VGND VPWR VPWR fd._0420_ sky130_fd_sc_hd__nand2_1
XFILLER_243_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_283_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4308_ fd._2496_ fd._2551_ fd._2562_ VGND VGND VPWR VPWR fd._2573_ sky130_fd_sc_hd__a21oi_1
XFILLER_82_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_1631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._8076_ fd._2423_ fd._2623_ fd._3398_ VGND VGND VPWR VPWR fd._3405_ sky130_fd_sc_hd__mux2_2
XFILLER_110_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5288_ fd._0082_ VGND VGND VPWR VPWR fd._0344_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_188_1691 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7027_ fd._1431_ fd._2255_ VGND VGND VPWR VPWR fd._2257_ sky130_fd_sc_hd__and2_1
Xfd._4239_ fd._1209_ fd.a\[3\] VGND VGND VPWR VPWR fd._1814_ sky130_fd_sc_hd__nor2b_1
XFILLER_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7929_ fd._3245_ fd._3248_ fd._3241_ VGND VGND VPWR VPWR fd._3249_ sky130_fd_sc_hd__mux2_1
XFILLER_109_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_278_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_269_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4590_ fd._3683_ fd._3535_ VGND VGND VPWR VPWR fd._3684_ sky130_fd_sc_hd__nor2_1
XFILLER_155_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_272_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_257_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6260_ fd._1405_ fd._1411_ fd._1412_ VGND VGND VPWR VPWR fd._1413_ sky130_fd_sc_hd__o21a_1
XFILLER_209_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_249_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5211_ fd._0256_ fd._0253_ fd._0255_ fd._0258_ VGND VGND VPWR VPWR fd._0259_ sky130_fd_sc_hd__a31oi_1
XFILLER_77_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6191_ fd._1329_ fd._1336_ VGND VGND VPWR VPWR fd._1337_ sky130_fd_sc_hd__and2_1
XTAP_4260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5142_ fd._4054_ fd._4061_ VGND VGND VPWR VPWR fd._0183_ sky130_fd_sc_hd__and2_1
XTAP_4293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5073_ fd._4005_ fd._4014_ VGND VGND VPWR VPWR fd._0107_ sky130_fd_sc_hd__or2b_1
XFILLER_162_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5975_ fd._0914_ fd._1098_ fd._1046_ VGND VGND VPWR VPWR fd._1100_ sky130_fd_sc_hd__mux2_1
XFILLER_186_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_277_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7714_ fd._2691_ fd._3011_ fd._2875_ VGND VGND VPWR VPWR fd._3012_ sky130_fd_sc_hd__mux2_1
Xfd._4926_ fd._3886_ fd._3858_ VGND VGND VPWR VPWR fd._4020_ sky130_fd_sc_hd__nand2_1
XFILLER_220_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_277_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_259_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._7645_ fd._2752_ fd._2757_ VGND VGND VPWR VPWR fd._2937_ sky130_fd_sc_hd__and2_1
XFILLER_133_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4857_ fd.b\[22\] fd._3949_ VGND VGND VPWR VPWR fd._3951_ sky130_fd_sc_hd__and2_1
XFILLER_173_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_250 VGND VGND VPWR VPWR user_project_wrapper_250/HI user_irq[0]
+ sky130_fd_sc_hd__conb_1
XFILLER_86_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_project_wrapper_261 VGND VGND VPWR VPWR user_project_wrapper_261/HI wbs_dat_o[7]
+ sky130_fd_sc_hd__conb_1
XFILLER_216_1518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_272 VGND VGND VPWR VPWR user_project_wrapper_272/HI wbs_dat_o[18]
+ sky130_fd_sc_hd__conb_1
XFILLER_82_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7576_ fd._2630_ fd._2860_ fd._2813_ VGND VGND VPWR VPWR fd._2861_ sky130_fd_sc_hd__mux2_1
Xuser_project_wrapper_283 VGND VGND VPWR VPWR user_project_wrapper_283/HI wbs_dat_o[29]
+ sky130_fd_sc_hd__conb_1
XFILLER_88_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4788_ fd._3675_ fd._3867_ VGND VGND VPWR VPWR fd._3882_ sky130_fd_sc_hd__nor2_1
XFILLER_173_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6527_ fd._1500_ fd._1706_ VGND VGND VPWR VPWR fd._1707_ sky130_fd_sc_hd__and2_1
XFILLER_141_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6458_ fd._1165_ fd._1630_ VGND VGND VPWR VPWR fd._1631_ sky130_fd_sc_hd__nand2_1
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5409_ fd._3947_ fd._0459_ VGND VGND VPWR VPWR fd._0477_ sky130_fd_sc_hd__nand2_1
XFILLER_283_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6389_ fd._1178_ fd._1554_ VGND VGND VPWR VPWR fd._1555_ sky130_fd_sc_hd__and2_1
XFILLER_244_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8128_ fd._3425_ fd._3434_ fd._3433_ VGND VGND VPWR VPWR fd._3443_ sky130_fd_sc_hd__a21o_1
XFILLER_270_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8059_ fd._3243_ fd._3256_ VGND VGND VPWR VPWR fd._3392_ sky130_fd_sc_hd__nand2_1
XFILLER_97_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_270_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_273_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_278_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_247_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_267_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5760_ fd._0862_ VGND VGND VPWR VPWR fd._0863_ sky130_fd_sc_hd__inv_2
XFILLER_7_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4711_ fd._3747_ fd._3645_ fd._3745_ VGND VGND VPWR VPWR fd._3805_ sky130_fd_sc_hd__and3_1
XFILLER_170_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5691_ fd._0782_ fd._0610_ VGND VGND VPWR VPWR fd._0787_ sky130_fd_sc_hd__xor2_1
XFILLER_100_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7430_ fd._2596_ fd._2699_ VGND VGND VPWR VPWR fd._2700_ sky130_fd_sc_hd__xnor2_1
Xfd._4642_ fd._3365_ fd._3735_ fd._3625_ VGND VGND VPWR VPWR fd._3736_ sky130_fd_sc_hd__mux2_1
XFILLER_135_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._7361_ fd._2426_ fd._2467_ VGND VGND VPWR VPWR fd._2624_ sky130_fd_sc_hd__nor2_1
XFILLER_257_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4573_ fd._3512_ fd._3666_ fd._3624_ VGND VGND VPWR VPWR fd._3667_ sky130_fd_sc_hd__mux2_1
XFILLER_215_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6312_ fd._0716_ fd._1468_ fd._1469_ VGND VGND VPWR VPWR fd._1470_ sky130_fd_sc_hd__a21oi_1
XFILLER_78_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7292_ fd._2547_ fd._2380_ VGND VGND VPWR VPWR fd._2548_ sky130_fd_sc_hd__and2_1
XFILLER_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6243_ fd._1211_ fd._1206_ VGND VGND VPWR VPWR fd._1394_ sky130_fd_sc_hd__or2_1
XFILLER_265_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_280_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6174_ fd._1062_ fd._1310_ fd._1073_ VGND VGND VPWR VPWR fd._1318_ sky130_fd_sc_hd__o21ai_1
XTAP_4090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5125_ fd._0156_ fd._0162_ fd._0163_ VGND VGND VPWR VPWR fd._0165_ sky130_fd_sc_hd__a21oi_1
XFILLER_94_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5056_ fd._3469_ VGND VGND VPWR VPWR fd._0089_ sky130_fd_sc_hd__buf_6
XFILLER_127_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_277_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5958_ fd._0933_ fd._1080_ VGND VGND VPWR VPWR fd._1081_ sky130_fd_sc_hd__xnor2_1
XFILLER_109_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_277_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._4909_ fd._4001_ fd._4002_ VGND VGND VPWR VPWR fd._4003_ sky130_fd_sc_hd__xnor2_1
XFILLER_175_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_256_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5889_ fd._0816_ fd._1004_ fd._0998_ VGND VGND VPWR VPWR fd._1005_ sky130_fd_sc_hd__mux2_1
XFILLER_133_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7628_ fd._1722_ fd._2917_ VGND VGND VPWR VPWR fd._2918_ sky130_fd_sc_hd__or2_1
XTAP_6409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7559_ fd._2840_ fd._2841_ VGND VGND VPWR VPWR fd._2842_ sky130_fd_sc_hd__nor2_1
XTAP_5719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_276_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_283_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_284_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_227_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_262_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_9035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_9046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_234_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_267_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6930_ fd._2141_ fd._2149_ VGND VGND VPWR VPWR fd._2150_ sky130_fd_sc_hd__and2_1
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6861_ fd._2055_ fd._2072_ VGND VGND VPWR VPWR fd._2074_ sky130_fd_sc_hd__or2_1
XFILLER_129_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5812_ fd._0684_ fd._0685_ VGND VGND VPWR VPWR fd._0920_ sky130_fd_sc_hd__and2_1
XFILLER_204_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_239_ fd.c\[31\] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_1
Xfd._6792_ fd._1729_ fd._1920_ fd._1785_ VGND VGND VPWR VPWR fd._1998_ sky130_fd_sc_hd__o21ai_1
XFILLER_200_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5743_ fd._0842_ fd._0799_ fd._0785_ VGND VGND VPWR VPWR fd._0844_ sky130_fd_sc_hd__o21a_1
XFILLER_170_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5674_ fd._0026_ VGND VGND VPWR VPWR fd._0768_ sky130_fd_sc_hd__buf_6
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_256_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_237_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7413_ fd._1286_ fd._2679_ VGND VGND VPWR VPWR fd._2681_ sky130_fd_sc_hd__or2_1
XFILLER_48_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4625_ fd._3625_ fd._3718_ VGND VGND VPWR VPWR fd._3719_ sky130_fd_sc_hd__nand2_1
XFILLER_174_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_1324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_258_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._7344_ fd._1666_ fd._2604_ VGND VGND VPWR VPWR fd._2605_ sky130_fd_sc_hd__and2_1
XFILLER_135_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._4556_ fd._3489_ fd._3649_ fd._3624_ VGND VGND VPWR VPWR fd._3650_ sky130_fd_sc_hd__mux2_1
XFILLER_170_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_284_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7275_ fd._2524_ fd._2528_ fd._2505_ VGND VGND VPWR VPWR fd._2530_ sky130_fd_sc_hd__mux2_1
XFILLER_284_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4487_ fd._3580_ fd._3233_ VGND VGND VPWR VPWR fd._3581_ sky130_fd_sc_hd__nand2_1
XFILLER_211_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6226_ fd._1372_ fd._1375_ fd._1349_ VGND VGND VPWR VPWR fd._1376_ sky130_fd_sc_hd__mux2_1
XFILLER_265_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_285_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_253_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6157_ fd._1148_ fd._1299_ VGND VGND VPWR VPWR fd._1300_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_263_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_253_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._5108_ fd._0088_ fd._0145_ VGND VGND VPWR VPWR fd._0146_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6088_ fd._0999_ fd._1222_ fd._1223_ VGND VGND VPWR VPWR fd._1224_ sky130_fd_sc_hd__mux2_1
XFILLER_181_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5039_ fd._1352_ fd._0069_ VGND VGND VPWR VPWR fd._0070_ sky130_fd_sc_hd__nand2_1
XFILLER_221_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_268_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_264_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_279_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_9 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_275_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_8164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4410_ fd._0252_ fd._1748_ VGND VGND VPWR VPWR fd._3504_ sky130_fd_sc_hd__or2_1
XTAP_7496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5390_ fd._0397_ fd._0402_ fd._0412_ VGND VGND VPWR VPWR fd._0456_ sky130_fd_sc_hd__a21o_1
XTAP_6773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._4341_ fd._1022_ fd._2837_ VGND VGND VPWR VPWR fd._2936_ sky130_fd_sc_hd__xnor2_1
XFILLER_208_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7060_ fd._2107_ fd._2292_ VGND VGND VPWR VPWR fd._2293_ sky130_fd_sc_hd__xor2_1
Xfd._4272_ fd._0197_ fd._2166_ VGND VGND VPWR VPWR fd._2177_ sky130_fd_sc_hd__xor2_1
XFILLER_212_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6011_ fd._1319_ fd._1137_ VGND VGND VPWR VPWR fd._1139_ sky130_fd_sc_hd__and2_1
XFILLER_63_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_267_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_263_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_85 VGND VGND VPWR VPWR user_project_wrapper_85/HI io_oeb[7]
+ sky130_fd_sc_hd__conb_1
XFILLER_21_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_96 VGND VGND VPWR VPWR user_project_wrapper_96/HI io_oeb[18]
+ sky130_fd_sc_hd__conb_1
XFILLER_235_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_250_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7962_ fd._3282_ fd._3284_ VGND VGND VPWR VPWR fd._3285_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_1659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6913_ fd._1722_ fd._2130_ VGND VGND VPWR VPWR fd._2131_ sky130_fd_sc_hd__nor2_1
XFILLER_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7893_ fd._0207_ fd._3085_ VGND VGND VPWR VPWR fd._3209_ sky130_fd_sc_hd__nor2_1
XFILLER_31_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6844_ fd._0965_ VGND VGND VPWR VPWR fd._2055_ sky130_fd_sc_hd__buf_6
XFILLER_239_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6775_ fd._0437_ fd._1821_ fd._1835_ fd._1915_ VGND VGND VPWR VPWR fd._1980_ sky130_fd_sc_hd__and4_1
XFILLER_239_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5726_ fd._0262_ fd._0825_ VGND VGND VPWR VPWR fd._0826_ sky130_fd_sc_hd__nand2_1
XFILLER_132_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_258_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5657_ fd._1264_ fd._0589_ VGND VGND VPWR VPWR fd._0750_ sky130_fd_sc_hd__and2_1
XFILLER_131_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_1356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4608_ fd._3671_ fd._3674_ fd._3701_ fd._3668_ VGND VGND VPWR VPWR fd._3702_ sky130_fd_sc_hd__o31a_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5588_ fd._0671_ fd._0672_ fd._0673_ VGND VGND VPWR VPWR fd._0674_ sky130_fd_sc_hd__or3_1
XFILLER_131_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_285_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_273_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7327_ fd._2332_ VGND VGND VPWR VPWR fd._2587_ sky130_fd_sc_hd__clkinv_2
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4539_ fd._3580_ fd._3632_ VGND VGND VPWR VPWR fd._3633_ sky130_fd_sc_hd__or2_1
XFILLER_245_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7258_ fd._2510_ fd._2393_ VGND VGND VPWR VPWR fd._2511_ sky130_fd_sc_hd__or2_1
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6209_ fd._1353_ fd._1356_ fd._1349_ VGND VGND VPWR VPWR fd._1357_ sky130_fd_sc_hd__mux2_1
XFILLER_25_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7189_ fd._2277_ fd._2275_ VGND VGND VPWR VPWR fd._2435_ sky130_fd_sc_hd__or2b_1
XFILLER_81_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput35 net35 VGND VGND VPWR VPWR io_out[10] sky130_fd_sc_hd__buf_2
XFILLER_150_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput46 net46 VGND VGND VPWR VPWR io_out[20] sky130_fd_sc_hd__buf_2
XFILLER_235_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput57 net57 VGND VGND VPWR VPWR io_out[30] sky130_fd_sc_hd__buf_2
XFILLER_27_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_277_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_264_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._4890_ fd._3868_ fd._3983_ fd._3882_ VGND VGND VPWR VPWR fd._3984_ sky130_fd_sc_hd__a21oi_1
XFILLER_201_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_279_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_275_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6560_ fd._1738_ fd._1742_ fd._1719_ VGND VGND VPWR VPWR fd._1743_ sky130_fd_sc_hd__mux2_1
XFILLER_99_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5511_ fd._0287_ fd._0588_ fd._0453_ VGND VGND VPWR VPWR fd._0589_ sky130_fd_sc_hd__mux2_1
XFILLER_154_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6491_ fd._1666_ fd._1664_ VGND VGND VPWR VPWR fd._1667_ sky130_fd_sc_hd__nor2_1
XFILLER_113_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._8230_ net70 net15 VGND VGND VPWR VPWR fd.a\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_239_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5442_ fd._0504_ fd._0511_ VGND VGND VPWR VPWR fd._0513_ sky130_fd_sc_hd__and2_1
XFILLER_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_282_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._8161_ fd._3475_ VGND VGND VPWR VPWR fd.ec\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_227_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5373_ fd._3689_ VGND VGND VPWR VPWR fd._0437_ sky130_fd_sc_hd__buf_6
XFILLER_132_1349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7112_ fd._2348_ fd._2349_ fd._2190_ VGND VGND VPWR VPWR fd._2350_ sky130_fd_sc_hd__a21bo_1
XFILLER_95_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_282_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4324_ fd._0010_ fd._1132_ VGND VGND VPWR VPWR fd._2749_ sky130_fd_sc_hd__nor2_1
XFILLER_212_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._8092_ fd._3414_ VGND VGND VPWR VPWR fd.mc\[13\] sky130_fd_sc_hd__clkbuf_1
XFILLER_94_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_282_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7043_ fd._2095_ fd._2272_ fd._2179_ fd._2273_ VGND VGND VPWR VPWR fd._2274_ sky130_fd_sc_hd__o31ai_2
XFILLER_251_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4255_ fd.b\[2\] fd._1924_ VGND VGND VPWR VPWR fd._1990_ sky130_fd_sc_hd__or2_1
XFILLER_47_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_251_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4186_ fd._1220_ VGND VGND VPWR VPWR fd._1231_ sky130_fd_sc_hd__buf_12
XFILLER_63_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7945_ fd._2377_ fd._1764_ fd._3265_ fd._2763_ VGND VGND VPWR VPWR fd._3267_ sky130_fd_sc_hd__a211o_1
XFILLER_91_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7876_ fd._2911_ VGND VGND VPWR VPWR fd._3191_ sky130_fd_sc_hd__clkinv_2
XFILLER_163_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6827_ fd._1242_ fd._2036_ VGND VGND VPWR VPWR fd._2037_ sky130_fd_sc_hd__nand2_1
XFILLER_50_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_258_1554 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._6758_ fd._1585_ fd._1771_ VGND VGND VPWR VPWR fd._1961_ sky130_fd_sc_hd__nor2_1
XFILLER_116_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_264_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_259_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5709_ fd._3883_ VGND VGND VPWR VPWR fd._0807_ sky130_fd_sc_hd__buf_6
XFILLER_172_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6689_ fd._1666_ fd._1868_ VGND VGND VPWR VPWR fd._1885_ sky130_fd_sc_hd__or2_1
XFILLER_132_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_269_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_259_1307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_259_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_276_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1663 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_264_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_281_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._5991_ fd._0716_ fd._1112_ fd._1116_ VGND VGND VPWR VPWR fd._1117_ sky130_fd_sc_hd__mux2_1
XFILLER_185_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4942_ fd._3853_ fd._3899_ VGND VGND VPWR VPWR fd._4036_ sky130_fd_sc_hd__nand2_1
XFILLER_220_1631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._7730_ fd._2481_ fd._2835_ VGND VGND VPWR VPWR fd._3030_ sky130_fd_sc_hd__nor2_1
XFILLER_9_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7661_ fd._2377_ fd._2765_ VGND VGND VPWR VPWR fd._2954_ sky130_fd_sc_hd__nand2_1
Xfd._4873_ fd._3773_ fd._3966_ VGND VGND VPWR VPWR fd._3967_ sky130_fd_sc_hd__and2_1
XFILLER_201_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6612_ fd._1798_ fd._1799_ VGND VGND VPWR VPWR fd._1800_ sky130_fd_sc_hd__nor2_1
Xfd._7592_ fd._2814_ fd._2877_ VGND VGND VPWR VPWR fd._2878_ sky130_fd_sc_hd__or2_1
XFILLER_114_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6543_ fd._0928_ fd._1546_ VGND VGND VPWR VPWR fd._1724_ sky130_fd_sc_hd__nor2_1
XFILLER_153_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_259_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6474_ fd._1464_ fd._1647_ fd._1615_ VGND VGND VPWR VPWR fd._1648_ sky130_fd_sc_hd__mux2_1
XFILLER_113_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_253_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8213_ net72 net28 VGND VGND VPWR VPWR fd.a\[5\] sky130_fd_sc_hd__dfxtp_1
Xfd._5425_ fd._0300_ fd._0493_ fd._0425_ VGND VGND VPWR VPWR fd._0495_ sky130_fd_sc_hd__mux2_1
XFILLER_214_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_283_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8144_ fd._3458_ VGND VGND VPWR VPWR fd.ec\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5356_ fd._0416_ fd._0418_ VGND VGND VPWR VPWR fd._0419_ sky130_fd_sc_hd__and2_1
XFILLER_95_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4307_ fd.b\[15\] fd._2540_ VGND VGND VPWR VPWR fd._2562_ sky130_fd_sc_hd__nor2_1
XFILLER_243_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8075_ fd._3403_ VGND VGND VPWR VPWR fd.mc\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_236_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5287_ fd._0868_ VGND VGND VPWR VPWR fd._0343_ sky130_fd_sc_hd__buf_6
XFILLER_184_1512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_247_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._7026_ fd._1431_ fd._2255_ VGND VGND VPWR VPWR fd._2256_ sky130_fd_sc_hd__nor2_1
XFILLER_63_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4238_ fd._0329_ fd._1781_ fd._1770_ fd._0307_ VGND VGND VPWR VPWR fd._1803_ sky130_fd_sc_hd__o211ai_1
XFILLER_208_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_251_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_260_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4169_ fd.b\[18\] fd._1033_ VGND VGND VPWR VPWR fd._1044_ sky130_fd_sc_hd__nor2_1
XFILLER_195_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7928_ fd._3246_ fd._3247_ VGND VGND VPWR VPWR fd._3248_ sky130_fd_sc_hd__xnor2_1
XFILLER_164_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7859_ fd._2876_ fd._3170_ fd._3165_ fd._3062_ fd._2763_ VGND VGND VPWR VPWR fd._3172_
+ sky130_fd_sc_hd__o221a_1
XFILLER_117_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_258_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_1663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_275_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_270_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_272_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_270_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5210_ fd._3689_ fd._0242_ fd._0244_ fd._4011_ VGND VGND VPWR VPWR fd._0258_ sky130_fd_sc_hd__a31oi_2
XFILLER_92_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6190_ fd._1334_ fd._1335_ VGND VGND VPWR VPWR fd._1336_ sky130_fd_sc_hd__nor2_1
XFILLER_77_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5141_ fd._0177_ fd._3646_ fd._0181_ VGND VGND VPWR VPWR fd._0182_ sky130_fd_sc_hd__mux2_1
XTAP_4283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5072_ fd._4010_ fd._4013_ VGND VGND VPWR VPWR fd._0106_ sky130_fd_sc_hd__or2_1
XFILLER_220_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_233_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5974_ fd._1097_ fd._0927_ VGND VGND VPWR VPWR fd._1098_ sky130_fd_sc_hd__xnor2_1
XFILLER_146_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7713_ fd._2806_ fd._3010_ VGND VGND VPWR VPWR fd._3011_ sky130_fd_sc_hd__xnor2_1
Xfd._4925_ fd._3990_ fd._3993_ fd._4018_ fd._3988_ VGND VGND VPWR VPWR fd._4019_ sky130_fd_sc_hd__o31a_1
XFILLER_146_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_255_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4856_ fd._3947_ fd._3949_ VGND VGND VPWR VPWR fd._3950_ sky130_fd_sc_hd__nor2_1
XFILLER_138_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7644_ fd._2933_ VGND VGND VPWR VPWR fd._2935_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_177_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_project_wrapper_240 VGND VGND VPWR VPWR user_project_wrapper_240/HI la_data_out[118]
+ sky130_fd_sc_hd__conb_1
XFILLER_255_1546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_251 VGND VGND VPWR VPWR user_project_wrapper_251/HI user_irq[1]
+ sky130_fd_sc_hd__conb_1
XFILLER_138_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_262 VGND VGND VPWR VPWR user_project_wrapper_262/HI wbs_dat_o[8]
+ sky130_fd_sc_hd__conb_1
XFILLER_245_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_273 VGND VGND VPWR VPWR user_project_wrapper_273/HI wbs_dat_o[19]
+ sky130_fd_sc_hd__conb_1
Xfd._4787_ fd._3869_ fd._3873_ fd._3879_ fd._3688_ fd._3880_ VGND VGND VPWR VPWR fd._3881_
+ sky130_fd_sc_hd__o221ai_2
Xfd._7575_ fd._2857_ fd._2858_ VGND VGND VPWR VPWR fd._2860_ sky130_fd_sc_hd__xnor2_1
Xuser_project_wrapper_284 VGND VGND VPWR VPWR user_project_wrapper_284/HI wbs_dat_o[30]
+ sky130_fd_sc_hd__conb_1
XFILLER_82_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6526_ fd._1498_ fd._1705_ VGND VGND VPWR VPWR fd._1706_ sky130_fd_sc_hd__nand2_1
XFILLER_29_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_275_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6457_ fd._1504_ fd._1629_ fd._1617_ VGND VGND VPWR VPWR fd._1630_ sky130_fd_sc_hd__mux2_1
XFILLER_60_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5408_ fd._0026_ fd._0475_ VGND VGND VPWR VPWR fd._0476_ sky130_fd_sc_hd__nor2_1
XFILLER_116_1697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6388_ fd._1548_ fd._1553_ fd._1533_ VGND VGND VPWR VPWR fd._1554_ sky130_fd_sc_hd__mux2_1
XFILLER_283_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8127_ fd._3440_ fd._3441_ VGND VGND VPWR VPWR fd._3442_ sky130_fd_sc_hd__nor2_1
XFILLER_244_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5339_ fd._0206_ fd._0399_ VGND VGND VPWR VPWR fd._0400_ sky130_fd_sc_hd__xnor2_1
XFILLER_82_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_266_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8058_ fd._3249_ fd._3388_ fd._3389_ fd._3390_ VGND VGND VPWR VPWR fd._3391_ sky130_fd_sc_hd__a22o_1
XFILLER_64_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_1304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7009_ fd._2236_ fd._2046_ VGND VGND VPWR VPWR fd._2237_ sky130_fd_sc_hd__xnor2_1
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_262_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_278_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_273_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_262_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout70 net71 VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_2
XFILLER_202_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4710_ fd._3645_ fd._3745_ fd._3747_ VGND VGND VPWR VPWR fd._3804_ sky130_fd_sc_hd__a21oi_1
XFILLER_143_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5690_ fd._3947_ VGND VGND VPWR VPWR fd._0786_ sky130_fd_sc_hd__buf_2
XFILLER_89_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_1522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4641_ fd._3640_ fd._3562_ VGND VGND VPWR VPWR fd._3735_ sky130_fd_sc_hd__xnor2_1
XFILLER_170_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7360_ fd._2506_ VGND VGND VPWR VPWR fd._2623_ sky130_fd_sc_hd__clkbuf_4
XFILLER_135_1528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4572_ fd._3664_ fd._3665_ VGND VGND VPWR VPWR fd._3666_ sky130_fd_sc_hd__xnor2_1
XFILLER_123_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_285_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_257_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6311_ fd._1448_ fd._1467_ VGND VGND VPWR VPWR fd._1469_ sky130_fd_sc_hd__nor2_1
XFILLER_2_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7291_ fd._1976_ fd._2545_ VGND VGND VPWR VPWR fd._2547_ sky130_fd_sc_hd__or2_1
XFILLER_215_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6242_ fd._3695_ fd._1392_ fd._1340_ fd._1348_ VGND VGND VPWR VPWR fd._1393_ sky130_fd_sc_hd__o211a_1
XFILLER_93_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6173_ fd._1051_ VGND VGND VPWR VPWR fd._1317_ sky130_fd_sc_hd__clkinv_2
XFILLER_64_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5124_ fd._3716_ fd._0161_ VGND VGND VPWR VPWR fd._0163_ sky130_fd_sc_hd__and2_1
XFILLER_209_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_280_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_252_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5055_ fd._3980_ fd._0086_ VGND VGND VPWR VPWR fd._0088_ sky130_fd_sc_hd__or2_1
XFILLER_166_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_1567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_277_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5957_ fd._0919_ fd._0925_ fd._0930_ VGND VGND VPWR VPWR fd._1080_ sky130_fd_sc_hd__o21a_1
XFILLER_107_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4908_ fd._3688_ fd._3879_ VGND VGND VPWR VPWR fd._4002_ sky130_fd_sc_hd__xnor2_1
XFILLER_238_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_277_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5888_ fd._0819_ fd._0836_ VGND VGND VPWR VPWR fd._1004_ sky130_fd_sc_hd__xnor2_1
XFILLER_259_1490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7627_ fd._2913_ fd._2916_ fd._2875_ VGND VGND VPWR VPWR fd._2917_ sky130_fd_sc_hd__mux2_1
XFILLER_133_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4839_ fd._3035_ fd._3794_ VGND VGND VPWR VPWR fd._3933_ sky130_fd_sc_hd__nand2_1
XFILLER_173_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_276_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7558_ fd._2657_ fd._2641_ fd._2656_ VGND VGND VPWR VPWR fd._2841_ sky130_fd_sc_hd__and3_1
XFILLER_138_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6509_ fd._1482_ fd._1686_ VGND VGND VPWR VPWR fd._1687_ sky130_fd_sc_hd__xnor2_1
XFILLER_134_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7489_ fd._1970_ fd._2670_ fd._2675_ VGND VGND VPWR VPWR fd._2765_ sky130_fd_sc_hd__and3_1
XFILLER_99_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_244_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_284_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_266_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_221_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_212_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_1601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_9058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_8357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_273_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_8379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_267_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_267_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_249_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6860_ fd._2055_ fd._2072_ VGND VGND VPWR VPWR fd._2073_ sky130_fd_sc_hd__nand2_1
XFILLER_204_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5811_ fd._0806_ fd._0810_ fd._0838_ fd._0804_ VGND VGND VPWR VPWR fd._0919_ sky130_fd_sc_hd__a31o_1
XFILLER_200_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_238_ fd.c\[30\] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6791_ fd._1986_ fd._1991_ fd._1993_ fd._1994_ fd._1996_ VGND VGND VPWR VPWR fd._1997_
+ sky130_fd_sc_hd__a2111o_1
XFILLER_278_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5742_ fd._0785_ fd._0842_ VGND VGND VPWR VPWR fd._0843_ sky130_fd_sc_hd__nor2_1
XFILLER_115_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_256_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_256_1641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5673_ fd._0026_ fd._0766_ VGND VGND VPWR VPWR fd._0767_ sky130_fd_sc_hd__or2_1
XFILLER_131_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4624_ fd._0857_ fd._3717_ VGND VGND VPWR VPWR fd._3718_ sky130_fd_sc_hd__xnor2_1
XFILLER_258_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_256_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7412_ fd._1286_ fd._2679_ VGND VGND VPWR VPWR fd._2680_ sky130_fd_sc_hd__nand2_1
XFILLER_174_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_258_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4555_ fd._3648_ fd._3546_ VGND VGND VPWR VPWR fd._3649_ sky130_fd_sc_hd__xor2_1
Xfd._7343_ fd._2409_ fd._2603_ fd._2506_ VGND VGND VPWR VPWR fd._2604_ sky130_fd_sc_hd__mux2_1
XFILLER_112_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_257_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7274_ fd._2525_ fd._2527_ VGND VGND VPWR VPWR fd._2528_ sky130_fd_sc_hd__xor2_1
XFILLER_272_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4486_ fd.b\[18\] VGND VGND VPWR VPWR fd._3580_ sky130_fd_sc_hd__buf_6
XFILLER_226_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_284_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6225_ fd._1196_ fd._1373_ VGND VGND VPWR VPWR fd._1375_ sky130_fd_sc_hd__xnor2_1
XFILLER_281_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6156_ fd._1155_ fd._1153_ VGND VGND VPWR VPWR fd._1299_ sky130_fd_sc_hd__or2b_1
XFILLER_65_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5107_ fd._3980_ fd._0086_ VGND VGND VPWR VPWR fd._0145_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6087_ fd._1169_ VGND VGND VPWR VPWR fd._1223_ sky130_fd_sc_hd__buf_6
XFILLER_263_1656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_1629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5038_ fd._0064_ fd._0066_ fd._0061_ fd._0068_ VGND VGND VPWR VPWR fd._0069_ sky130_fd_sc_hd__a31o_1
XFILLER_181_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_267_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6989_ fd._1933_ fd._1997_ fd._2214_ VGND VGND VPWR VPWR fd._2215_ sky130_fd_sc_hd__and3_1
XFILLER_162_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_270_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_263_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_240_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_275_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4340_ fd.b\[19\] fd._2914_ VGND VGND VPWR VPWR fd._2925_ sky130_fd_sc_hd__and2_1
XTAP_6796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4271_ fd._0186_ fd._2089_ fd._1341_ fd.a\[6\] VGND VGND VPWR VPWR fd._2166_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_169_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_281_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_267_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6010_ fd._1308_ fd._1137_ VGND VGND VPWR VPWR fd._1138_ sky130_fd_sc_hd__or2_1
XFILLER_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_project_wrapper_86 VGND VGND VPWR VPWR user_project_wrapper_86/HI io_oeb[8]
+ sky130_fd_sc_hd__conb_1
XFILLER_62_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_97 VGND VGND VPWR VPWR user_project_wrapper_97/HI io_oeb[19]
+ sky130_fd_sc_hd__conb_1
XFILLER_37_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_250_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7961_ fd._3283_ fd._3163_ VGND VGND VPWR VPWR fd._3284_ sky130_fd_sc_hd__nand2_1
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6912_ fd._2129_ VGND VGND VPWR VPWR fd._2130_ sky130_fd_sc_hd__inv_2
XFILLER_124_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7892_ fd._1286_ fd._3092_ VGND VGND VPWR VPWR fd._3208_ sky130_fd_sc_hd__and2_1
XFILLER_15_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6843_ fd._0131_ fd._2053_ VGND VGND VPWR VPWR fd._2054_ sky130_fd_sc_hd__nor2_1
XFILLER_198_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6774_ fd._1821_ fd._1835_ fd._1915_ fd._1977_ VGND VGND VPWR VPWR fd._1978_ sky130_fd_sc_hd__a31o_1
XFILLER_274_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5725_ fd._0636_ fd._0823_ fd._0801_ VGND VGND VPWR VPWR fd._0825_ sky130_fd_sc_hd__mux2_1
XFILLER_171_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5656_ fd._0000_ fd._0744_ fd._0746_ fd._0748_ VGND VGND VPWR VPWR fd._0749_ sky130_fd_sc_hd__a211o_1
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_258_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._4607_ fd._3682_ fd._3699_ fd._3700_ fd._3680_ VGND VGND VPWR VPWR fd._3701_ sky130_fd_sc_hd__o211a_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5587_ fd._0521_ fd._0524_ fd._0514_ VGND VGND VPWR VPWR fd._0673_ sky130_fd_sc_hd__a21oi_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7326_ fd._1102_ fd._2585_ fd._2582_ fd._2576_ VGND VGND VPWR VPWR fd._2586_ sky130_fd_sc_hd__o2bb2a_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4538_ fd._3571_ fd._3631_ fd._3625_ VGND VGND VPWR VPWR fd._3632_ sky130_fd_sc_hd__mux2_1
XFILLER_257_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4469_ fd._3449_ fd._3560_ fd._3562_ fd._3430_ VGND VGND VPWR VPWR fd._3563_ sky130_fd_sc_hd__or4_1
XFILLER_211_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7257_ fd._2395_ VGND VGND VPWR VPWR fd._2510_ sky130_fd_sc_hd__clkinv_2
XFILLER_72_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_285_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6208_ fd._1218_ fd._1355_ VGND VGND VPWR VPWR fd._1356_ sky130_fd_sc_hd__xnor2_1
XFILLER_26_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_281_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7188_ fd._2427_ fd._2433_ VGND VGND VPWR VPWR fd._2434_ sky130_fd_sc_hd__nand2_1
XFILLER_25_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_285_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6139_ fd._1115_ fd._1279_ fd._1223_ VGND VGND VPWR VPWR fd._1280_ sky130_fd_sc_hd__mux2_1
XFILLER_20_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_257_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput36 net36 VGND VGND VPWR VPWR io_out[11] sky130_fd_sc_hd__buf_2
XFILLER_134_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput47 net47 VGND VGND VPWR VPWR io_out[21] sky130_fd_sc_hd__buf_2
XFILLER_235_1533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput58 net58 VGND VGND VPWR VPWR io_out[31] sky130_fd_sc_hd__buf_2
XFILLER_0_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_1515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_1559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_1368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5510_ fd._0587_ VGND VGND VPWR VPWR fd._0588_ sky130_fd_sc_hd__clkinv_2
XFILLER_153_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6490_ fd._0758_ VGND VGND VPWR VPWR fd._1666_ sky130_fd_sc_hd__buf_6
XTAP_7250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_1628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5441_ fd._0504_ fd._0511_ VGND VGND VPWR VPWR fd._0512_ sky130_fd_sc_hd__nor2_1
XFILLER_136_1464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_1639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5372_ fd._0262_ fd._0435_ VGND VGND VPWR VPWR fd._0436_ sky130_fd_sc_hd__nand2_1
Xfd._8160_ fd._3473_ fd._3474_ VGND VGND VPWR VPWR fd._3475_ sky130_fd_sc_hd__or2_1
XFILLER_239_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_282_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4323_ fd._4049_ VGND VGND VPWR VPWR fd._2738_ sky130_fd_sc_hd__buf_6
XTAP_5881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7111_ fd._2174_ fd._2189_ VGND VGND VPWR VPWR fd._2349_ sky130_fd_sc_hd__nor2_1
XTAP_5892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._8091_ fd._1047_ fd._1232_ fd._3411_ VGND VGND VPWR VPWR fd._3414_ sky130_fd_sc_hd__mux2_1
XFILLER_54_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4254_ fd.b\[1\] fd._1946_ fd._1957_ VGND VGND VPWR VPWR fd._1979_ sky130_fd_sc_hd__or3_1
XFILLER_184_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._7042_ fd._2090_ fd._2179_ VGND VGND VPWR VPWR fd._2273_ sky130_fd_sc_hd__nand2_1
XFILLER_263_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_282_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_251_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4185_ fd._1209_ VGND VGND VPWR VPWR fd._1220_ sky130_fd_sc_hd__buf_8
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7944_ fd._1764_ fd._3077_ VGND VGND VPWR VPWR fd._3265_ sky130_fd_sc_hd__nor2_1
XFILLER_17_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7875_ fd._3136_ fd._3140_ fd._3180_ fd._3187_ fd._3188_ VGND VGND VPWR VPWR fd._3190_
+ sky130_fd_sc_hd__o41a_1
XFILLER_191_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6826_ fd._1828_ fd._2035_ fd._2020_ VGND VGND VPWR VPWR fd._2036_ sky130_fd_sc_hd__mux2_1
XFILLER_144_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._6757_ fd._1397_ fd._1959_ VGND VGND VPWR VPWR fd._1960_ sky130_fd_sc_hd__nand2_1
XFILLER_171_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5708_ fd._0804_ fd._0805_ VGND VGND VPWR VPWR fd._0806_ sky130_fd_sc_hd__nor2_1
XFILLER_67_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6688_ fd._1796_ fd._1799_ fd._1882_ fd._1883_ VGND VGND VPWR VPWR fd._1884_ sky130_fd_sc_hd__o211ai_2
XFILLER_259_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5639_ fd._4055_ fd._0729_ VGND VGND VPWR VPWR fd._0730_ sky130_fd_sc_hd__xnor2_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7309_ fd._2344_ VGND VGND VPWR VPWR fd._2567_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_280_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_259_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_276_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_276_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5990_ fd._1451_ fd._1115_ VGND VGND VPWR VPWR fd._1116_ sky130_fd_sc_hd__xnor2_1
XFILLER_158_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4941_ fd._3982_ fd._4028_ fd._4033_ fd._4034_ VGND VGND VPWR VPWR fd._4035_ sky130_fd_sc_hd__a31o_1
XFILLER_201_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7660_ fd._1970_ fd._2813_ VGND VGND VPWR VPWR fd._2953_ sky130_fd_sc_hd__nand2_1
Xfd._4872_ fd._3794_ fd._3965_ fd._3960_ VGND VGND VPWR VPWR fd._3966_ sky130_fd_sc_hd__mux2_1
XFILLER_220_1676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6611_ fd._1797_ fd._1721_ VGND VGND VPWR VPWR fd._1799_ sky130_fd_sc_hd__nor2_1
XFILLER_160_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7591_ fd._2875_ VGND VGND VPWR VPWR fd._2877_ sky130_fd_sc_hd__buf_6
XFILLER_173_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6542_ fd._1558_ fd._1566_ fd._1596_ fd._1555_ VGND VGND VPWR VPWR fd._1723_ sky130_fd_sc_hd__a31o_1
XFILLER_64_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._6473_ fd._1459_ fd._1646_ VGND VGND VPWR VPWR fd._1647_ sky130_fd_sc_hd__xnor2_1
XFILLER_45_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8212_ net72 net27 VGND VGND VPWR VPWR fd.a\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_256_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5424_ fd._0341_ fd._0485_ VGND VGND VPWR VPWR fd._0493_ sky130_fd_sc_hd__xnor2_1
XFILLER_45_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_282_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8143_ fd._3456_ fd._3457_ VGND VGND VPWR VPWR fd._3458_ sky130_fd_sc_hd__or2_1
XFILLER_94_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5355_ fd._3773_ fd._0415_ VGND VGND VPWR VPWR fd._0418_ sky130_fd_sc_hd__or2_1
XFILLER_209_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_1600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_282_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4306_ fd.b\[15\] fd._2540_ VGND VGND VPWR VPWR fd._2551_ sky130_fd_sc_hd__nand2_1
XFILLER_247_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5286_ fd._0330_ fd._0336_ fd._0337_ fd._0338_ fd._0341_ VGND VGND VPWR VPWR fd._0342_
+ sky130_fd_sc_hd__a2111o_1
Xfd._8074_ fd._2623_ fd._2813_ fd._3398_ VGND VGND VPWR VPWR fd._3403_ sky130_fd_sc_hd__mux2_2
XFILLER_188_1671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7025_ fd._2065_ fd._2253_ fd._2116_ VGND VGND VPWR VPWR fd._2255_ sky130_fd_sc_hd__mux2_1
XFILLER_251_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4237_ fd._0307_ fd._1770_ fd._1781_ fd._0329_ VGND VGND VPWR VPWR fd._1792_ sky130_fd_sc_hd__a211o_1
XFILLER_282_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._4168_ fd.a\[18\] VGND VGND VPWR VPWR fd._1033_ sky130_fd_sc_hd__inv_2
XFILLER_251_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4099_ fd._0241_ fd._0263_ VGND VGND VPWR VPWR fd._0274_ sky130_fd_sc_hd__nor2_1
XFILLER_91_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7927_ fd._3228_ fd._3221_ VGND VGND VPWR VPWR fd._3247_ sky130_fd_sc_hd__and2b_1
XFILLER_143_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7858_ fd._1211_ fd._3170_ VGND VGND VPWR VPWR fd._3171_ sky130_fd_sc_hd__nand2_1
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6809_ fd._2016_ fd._1910_ fd._1829_ VGND VGND VPWR VPWR fd._2017_ sky130_fd_sc_hd__o21a_1
XFILLER_117_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7789_ fd._3005_ fd._3094_ fd._3076_ VGND VGND VPWR VPWR fd._3095_ sky130_fd_sc_hd__mux2_1
XFILLER_145_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_259_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1670 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_262_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_1676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_278_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_276_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_264_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5140_ fd._4055_ fd._0180_ VGND VGND VPWR VPWR fd._0181_ sky130_fd_sc_hd__xnor2_1
XFILLER_168_1519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5071_ fd._0104_ VGND VGND VPWR VPWR fd._0105_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_217_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5973_ fd._0933_ fd._1080_ fd._0909_ VGND VGND VPWR VPWR fd._1097_ sky130_fd_sc_hd__a21o_1
XFILLER_185_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7712_ fd._2698_ fd._2803_ VGND VGND VPWR VPWR fd._3010_ sky130_fd_sc_hd__nand2_1
XFILLER_9_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4924_ fd._3999_ fd._4015_ fd._4016_ fd._4017_ VGND VGND VPWR VPWR fd._4018_ sky130_fd_sc_hd__o211a_1
XFILLER_179_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7643_ fd._2533_ fd._2933_ VGND VGND VPWR VPWR fd._2934_ sky130_fd_sc_hd__nand2_1
Xfd._4855_ fd._3776_ fd._3948_ fd._3800_ VGND VGND VPWR VPWR fd._3949_ sky130_fd_sc_hd__mux2_1
XFILLER_161_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_230 VGND VGND VPWR VPWR user_project_wrapper_230/HI la_data_out[108]
+ sky130_fd_sc_hd__conb_1
XFILLER_154_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_project_wrapper_241 VGND VGND VPWR VPWR user_project_wrapper_241/HI la_data_out[119]
+ sky130_fd_sc_hd__conb_1
Xuser_project_wrapper_252 VGND VGND VPWR VPWR user_project_wrapper_252/HI user_irq[2]
+ sky130_fd_sc_hd__conb_1
XFILLER_160_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7574_ fd._1507_ fd._2627_ VGND VGND VPWR VPWR fd._2858_ sky130_fd_sc_hd__xnor2_1
XFILLER_138_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_project_wrapper_263 VGND VGND VPWR VPWR user_project_wrapper_263/HI wbs_dat_o[9]
+ sky130_fd_sc_hd__conb_1
XFILLER_255_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._4786_ fd._3688_ fd._3878_ fd._3875_ fd.b\[1\] VGND VGND VPWR VPWR fd._3880_ sky130_fd_sc_hd__a211o_1
XFILLER_114_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_274 VGND VGND VPWR VPWR user_project_wrapper_274/HI wbs_dat_o[20]
+ sky130_fd_sc_hd__conb_1
XFILLER_245_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_285 VGND VGND VPWR VPWR user_project_wrapper_285/HI wbs_dat_o[31]
+ sky130_fd_sc_hd__conb_1
Xfd._6525_ fd._1438_ fd._1496_ fd._1499_ VGND VGND VPWR VPWR fd._1705_ sky130_fd_sc_hd__a21o_1
XFILLER_173_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6456_ fd._1425_ fd._1628_ VGND VGND VPWR VPWR fd._1629_ sky130_fd_sc_hd__xor2_1
XFILLER_151_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_256_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5407_ fd._0400_ fd._0474_ fd._0453_ VGND VGND VPWR VPWR fd._0475_ sky130_fd_sc_hd__mux2_1
XFILLER_151_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_283_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6387_ fd._1549_ fd._1552_ VGND VGND VPWR VPWR fd._1553_ sky130_fd_sc_hd__xor2_1
XFILLER_99_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_1580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8126_ fd.a\[25\] fd.b\[25\] VGND VGND VPWR VPWR fd._3441_ sky130_fd_sc_hd__and2b_1
XFILLER_55_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5338_ fd._0242_ fd._0244_ fd._0398_ VGND VGND VPWR VPWR fd._0399_ sky130_fd_sc_hd__a21oi_1
XFILLER_209_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_1632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8057_ fd._3221_ fd._3230_ fd._3235_ VGND VGND VPWR VPWR fd._3390_ sky130_fd_sc_hd__nand3_1
XFILLER_24_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5269_ fd._0118_ fd._0322_ fd._0268_ VGND VGND VPWR VPWR fd._0323_ sky130_fd_sc_hd__mux2_1
XFILLER_3_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7008_ fd._2037_ fd._2235_ fd._2043_ VGND VGND VPWR VPWR fd._2236_ sky130_fd_sc_hd__a21o_1
XFILLER_145_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_8528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_262_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_261_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout71 net75 VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__buf_2
XFILLER_230_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4640_ fd._3646_ VGND VGND VPWR VPWR fd._3734_ sky130_fd_sc_hd__clkinv_4
XFILLER_142_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_252_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_269_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4571_ fd._3513_ fd._3542_ VGND VGND VPWR VPWR fd._3665_ sky130_fd_sc_hd__nand2_1
XFILLER_69_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6310_ fd._1448_ fd._1467_ VGND VGND VPWR VPWR fd._1468_ sky130_fd_sc_hd__xor2_1
XFILLER_46_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7290_ fd._2545_ VGND VGND VPWR VPWR fd._2546_ sky130_fd_sc_hd__clkinv_2
XFILLER_111_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_265_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6241_ fd._1232_ VGND VGND VPWR VPWR fd._1392_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_42_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6172_ fd._1314_ fd._1315_ VGND VGND VPWR VPWR fd._1316_ sky130_fd_sc_hd__nand2_1
XTAP_4070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5123_ fd._3716_ fd._0161_ VGND VGND VPWR VPWR fd._0162_ sky130_fd_sc_hd__or2_1
XFILLER_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_283_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5054_ fd._0085_ fd._4023_ fd._0060_ VGND VGND VPWR VPWR fd._0086_ sky130_fd_sc_hd__mux2_1
XFILLER_166_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_1669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_1579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_1412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5956_ fd._1075_ fd._1062_ fd._1078_ VGND VGND VPWR VPWR fd._1079_ sky130_fd_sc_hd__or3_1
XFILLER_88_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_277_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4907_ fd.b\[1\] fd._3875_ VGND VGND VPWR VPWR fd._4001_ sky130_fd_sc_hd__or2_1
XFILLER_106_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5887_ fd._1001_ fd._1002_ VGND VGND VPWR VPWR fd._1003_ sky130_fd_sc_hd__nand2_1
XFILLER_162_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7626_ fd._2773_ fd._2915_ VGND VGND VPWR VPWR fd._2916_ sky130_fd_sc_hd__xnor2_1
Xfd._4838_ fd._3808_ fd._3930_ fd._3931_ VGND VGND VPWR VPWR fd._3932_ sky130_fd_sc_hd__or3_1
XFILLER_115_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7557_ fd._2641_ fd._2656_ fd._2657_ VGND VGND VPWR VPWR fd._2840_ sky130_fd_sc_hd__a21oi_1
Xfd._4769_ fd._3694_ fd._3697_ VGND VGND VPWR VPWR fd._3863_ sky130_fd_sc_hd__and2_1
XFILLER_170_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_275_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6508_ fd._1492_ fd._1488_ VGND VGND VPWR VPWR fd._1686_ sky130_fd_sc_hd__and2b_1
XFILLER_29_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_272_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7488_ fd._2759_ fd._2762_ fd._2763_ VGND VGND VPWR VPWR fd._2764_ sky130_fd_sc_hd__o21a_1
XFILLER_275_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6439_ fd._1102_ fd._1535_ VGND VGND VPWR VPWR fd._1610_ sky130_fd_sc_hd__nor2_1
XFILLER_112_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8109_ fd._3621_ fd._3626_ fd._3222_ VGND VGND VPWR VPWR fd.mc\[22\] sky130_fd_sc_hd__o21a_1
XFILLER_244_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_243_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_266_1495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_221_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_245_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_260_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_1668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_278_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_1636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5810_ fd._0910_ fd._0915_ fd._0917_ VGND VGND VPWR VPWR fd._0918_ sky130_fd_sc_hd__a21o_1
X_237_ fd.c\[29\] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_1
XFILLER_15_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6790_ fd._1931_ fd._1995_ VGND VGND VPWR VPWR fd._1996_ sky130_fd_sc_hd__nand2_1
XFILLER_128_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5741_ fd._0841_ fd._0792_ fd._0790_ VGND VGND VPWR VPWR fd._0842_ sky130_fd_sc_hd__o21a_1
XFILLER_183_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5672_ fd._0605_ fd._0765_ VGND VGND VPWR VPWR fd._0766_ sky130_fd_sc_hd__xnor2_1
XFILLER_170_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7411_ fd._2622_ fd._2677_ fd._2678_ VGND VGND VPWR VPWR fd._2679_ sky130_fd_sc_hd__a21oi_2
XTAP_8881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4623_ fd._3498_ fd._3549_ VGND VGND VPWR VPWR fd._3717_ sky130_fd_sc_hd__nand2_1
XFILLER_217_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7342_ fd._2404_ fd._2602_ VGND VGND VPWR VPWR fd._2603_ sky130_fd_sc_hd__xnor2_1
XFILLER_26_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4554_ fd._3548_ fd._3647_ fd._3496_ VGND VGND VPWR VPWR fd._3648_ sky130_fd_sc_hd__o21ai_1
XFILLER_65_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_273_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7273_ fd._2526_ fd._2385_ VGND VGND VPWR VPWR fd._2527_ sky130_fd_sc_hd__nor2_1
XFILLER_38_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4485_ fd.b\[18\] fd._3233_ VGND VGND VPWR VPWR fd._3579_ sky130_fd_sc_hd__or2_1
XFILLER_61_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6224_ fd._1205_ fd._1213_ VGND VGND VPWR VPWR fd._1373_ sky130_fd_sc_hd__and2_1
XFILLER_93_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_265_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_281_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6155_ fd._1233_ fd._1295_ fd._1296_ VGND VGND VPWR VPWR fd._1298_ sky130_fd_sc_hd__a21oi_1
XFILLER_20_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_280_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5106_ fd._3708_ fd._0139_ VGND VGND VPWR VPWR fd._0144_ sky130_fd_sc_hd__nand2_1
XFILLER_209_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6086_ fd._1034_ fd._1221_ VGND VGND VPWR VPWR fd._1222_ sky130_fd_sc_hd__nand2_1
XFILLER_185_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5037_ fd._0013_ fd._0067_ VGND VGND VPWR VPWR fd._0068_ sky130_fd_sc_hd__and2_1
XFILLER_221_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_261_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6988_ fd._2004_ fd._2003_ VGND VGND VPWR VPWR fd._2214_ sky130_fd_sc_hd__or2b_1
XFILLER_179_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5939_ fd._1040_ fd._0981_ VGND VGND VPWR VPWR fd._1060_ sky130_fd_sc_hd__xnor2_1
XFILLER_88_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_283_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7609_ fd._2712_ fd._2794_ VGND VGND VPWR VPWR fd._2897_ sky130_fd_sc_hd__xnor2_1
XTAP_6219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_276_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_1568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_279_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4270_ fd.b\[8\] VGND VGND VPWR VPWR fd._2155_ sky130_fd_sc_hd__buf_6
XFILLER_212_1578 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_281_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_263_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_project_wrapper_87 VGND VGND VPWR VPWR user_project_wrapper_87/HI io_oeb[9]
+ sky130_fd_sc_hd__conb_1
XFILLER_165_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_project_wrapper_98 VGND VGND VPWR VPWR user_project_wrapper_98/HI io_oeb[20]
+ sky130_fd_sc_hd__conb_1
XFILLER_267_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7960_ fd._2751_ fd._3162_ VGND VGND VPWR VPWR fd._3283_ sky130_fd_sc_hd__nand2_1
XFILLER_15_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_1376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_231_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6911_ fd._1989_ fd._2128_ fd._2115_ VGND VGND VPWR VPWR fd._2129_ sky130_fd_sc_hd__mux2_1
XFILLER_128_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7891_ fd._3105_ fd._3122_ fd._3203_ fd._3206_ VGND VGND VPWR VPWR fd._3207_ sky130_fd_sc_hd__a31o_1
XFILLER_31_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6842_ fd._2052_ VGND VGND VPWR VPWR fd._2053_ sky130_fd_sc_hd__inv_2
XFILLER_89_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_274_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6773_ fd._1961_ fd._1972_ VGND VGND VPWR VPWR fd._1977_ sky130_fd_sc_hd__or2b_1
XFILLER_7_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5724_ fd._0820_ fd._0822_ VGND VGND VPWR VPWR fd._0823_ sky130_fd_sc_hd__xor2_1
XFILLER_144_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5655_ fd._0739_ fd._0742_ VGND VGND VPWR VPWR fd._0748_ sky130_fd_sc_hd__and2_1
XFILLER_135_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4606_ fd._0252_ fd._3673_ VGND VGND VPWR VPWR fd._3700_ sky130_fd_sc_hd__or2_1
XFILLER_112_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5586_ fd._0465_ fd._0481_ fd._0612_ VGND VGND VPWR VPWR fd._0672_ sky130_fd_sc_hd__and3_2
XFILLER_285_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7325_ fd._2576_ fd._2583_ VGND VGND VPWR VPWR fd._2585_ sky130_fd_sc_hd__xnor2_1
XFILLER_131_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4537_ fd._3630_ fd._3573_ VGND VGND VPWR VPWR fd._3631_ sky130_fd_sc_hd__xnor2_1
XFILLER_135_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._7256_ fd._1330_ fd._2508_ VGND VGND VPWR VPWR fd._2509_ sky130_fd_sc_hd__or2_1
XFILLER_2_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4468_ fd._3376_ fd._3561_ VGND VGND VPWR VPWR fd._3562_ sky130_fd_sc_hd__nand2_1
XFILLER_6_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6207_ fd._1226_ fd._1354_ VGND VGND VPWR VPWR fd._1355_ sky130_fd_sc_hd__nand2_1
XFILLER_96_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_285_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7187_ fd._2260_ fd._2432_ fd._2323_ VGND VGND VPWR VPWR fd._2433_ sky130_fd_sc_hd__mux2_1
Xfd._4399_ fd._3492_ fd._2122_ VGND VGND VPWR VPWR fd._3493_ sky130_fd_sc_hd__nor2_1
XFILLER_241_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_281_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6138_ fd._1112_ fd._1116_ VGND VGND VPWR VPWR fd._1279_ sky130_fd_sc_hd__xor2_1
XFILLER_228_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6069_ fd._1200_ fd._1202_ VGND VGND VPWR VPWR fd._1203_ sky130_fd_sc_hd__xnor2_1
XFILLER_224_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_257_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput37 net37 VGND VGND VPWR VPWR io_out[12] sky130_fd_sc_hd__buf_2
XFILLER_162_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_270_1403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput48 net48 VGND VGND VPWR VPWR io_out[22] sky130_fd_sc_hd__buf_2
XFILLER_153_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_270_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_1545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput59 net59 VGND VGND VPWR VPWR io_out[3] sky130_fd_sc_hd__buf_2
XFILLER_235_1556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_277_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_263_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_1663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_1527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_253_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_1656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5440_ fd._0506_ fd._0510_ fd._0425_ VGND VGND VPWR VPWR fd._0511_ sky130_fd_sc_hd__mux2_1
XFILLER_239_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5371_ fd._0431_ fd._0434_ fd._0425_ VGND VGND VPWR VPWR fd._0435_ sky130_fd_sc_hd__mux2_1
XTAP_6583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7110_ fd._2142_ fd._2164_ VGND VGND VPWR VPWR fd._2348_ sky130_fd_sc_hd__or2_1
Xfd._4322_ fd._2672_ fd._2716_ VGND VGND VPWR VPWR fd._2727_ sky130_fd_sc_hd__xnor2_1
XFILLER_94_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8090_ fd._3413_ VGND VGND VPWR VPWR fd.mc\[12\] sky130_fd_sc_hd__clkbuf_1
XFILLER_212_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7041_ fd._2271_ fd._2092_ VGND VGND VPWR VPWR fd._2272_ sky130_fd_sc_hd__nor2_1
Xfd._4253_ fd._1946_ fd._1957_ fd.b\[1\] VGND VGND VPWR VPWR fd._1968_ sky130_fd_sc_hd__o21a_1
XFILLER_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4184_ fd._4060_ fd._1187_ fd._1198_ VGND VGND VPWR VPWR fd._1209_ sky130_fd_sc_hd__a21o_4
XFILLER_63_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_250_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_250_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7943_ fd._3243_ fd._3256_ fd._3262_ fd._3263_ VGND VGND VPWR VPWR fd._3264_ sky130_fd_sc_hd__and4_1
XFILLER_203_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7874_ fd._3185_ fd._3132_ fd._3184_ VGND VGND VPWR VPWR fd._3188_ sky130_fd_sc_hd__o21bai_1
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6825_ fd._2016_ fd._1911_ VGND VGND VPWR VPWR fd._2035_ sky130_fd_sc_hd__xnor2_1
XFILLER_129_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6756_ fd._1813_ fd._1763_ fd._1766_ VGND VGND VPWR VPWR fd._1959_ sky130_fd_sc_hd__o21ai_1
XFILLER_116_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5707_ fd._1341_ fd._0803_ VGND VGND VPWR VPWR fd._0805_ sky130_fd_sc_hd__nor2_1
XFILLER_171_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6687_ fd._1798_ VGND VGND VPWR VPWR fd._1883_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_154_1510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_259_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5638_ fd._0562_ fd._0728_ fd._0614_ VGND VGND VPWR VPWR fd._0729_ sky130_fd_sc_hd__mux2_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_258_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5569_ fd._1264_ fd._0652_ VGND VGND VPWR VPWR fd._0653_ sky130_fd_sc_hd__or2_1
XFILLER_140_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_285_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7308_ fd._1600_ VGND VGND VPWR VPWR fd._2566_ sky130_fd_sc_hd__clkbuf_2
XFILLER_6_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_261_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7239_ fd._2297_ fd._2304_ VGND VGND VPWR VPWR fd._2490_ sky130_fd_sc_hd__xnor2_1
XFILLER_26_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_257_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_272_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_283_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4940_ fd._0868_ fd._4032_ VGND VGND VPWR VPWR fd._4034_ sky130_fd_sc_hd__nor2_1
XFILLER_125_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4871_ fd._3935_ fd._3964_ VGND VGND VPWR VPWR fd._3965_ sky130_fd_sc_hd__nand2_1
XFILLER_8_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6610_ fd._1797_ fd._1721_ VGND VGND VPWR VPWR fd._1798_ sky130_fd_sc_hd__and2_1
XFILLER_275_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7590_ fd._2875_ VGND VGND VPWR VPWR fd._2876_ sky130_fd_sc_hd__clkinv_8
XFILLER_99_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_275_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6541_ fd._0662_ VGND VGND VPWR VPWR fd._1722_ sky130_fd_sc_hd__buf_6
XFILLER_153_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_253_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_1598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6472_ fd._1466_ fd._1465_ VGND VGND VPWR VPWR fd._1646_ sky130_fd_sc_hd__and2b_1
XTAP_7070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8211_ net72 net26 VGND VGND VPWR VPWR fd.a\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_7092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5423_ fd._0489_ fd._0491_ VGND VGND VPWR VPWR fd._0492_ sky130_fd_sc_hd__nor2_1
XFILLER_136_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8142_ fd._3447_ fd._3455_ VGND VGND VPWR VPWR fd._3457_ sky130_fd_sc_hd__and2_1
Xfd._5354_ fd._3773_ fd._0415_ VGND VGND VPWR VPWR fd._0416_ sky130_fd_sc_hd__nand2_1
XFILLER_7_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_255_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_282_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4305_ fd._2507_ fd._2529_ fd._1231_ VGND VGND VPWR VPWR fd._2540_ sky130_fd_sc_hd__mux2_1
XFILLER_3_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8073_ fd._3402_ VGND VGND VPWR VPWR fd.mc\[4\] sky130_fd_sc_hd__clkbuf_1
XFILLER_282_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5285_ fd._0301_ fd._0339_ VGND VGND VPWR VPWR fd._0341_ sky130_fd_sc_hd__nand2_1
XFILLER_264_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7024_ fd._2251_ fd._2252_ VGND VGND VPWR VPWR fd._2253_ sky130_fd_sc_hd__xnor2_1
XFILLER_63_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4236_ fd._0351_ fd._0395_ VGND VGND VPWR VPWR fd._1781_ sky130_fd_sc_hd__and2_1
XFILLER_24_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._4167_ fd._0032_ fd._0109_ VGND VGND VPWR VPWR fd._1022_ sky130_fd_sc_hd__or2_1
XFILLER_260_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4098_ fd._0252_ fd.a\[5\] VGND VGND VPWR VPWR fd._0263_ sky130_fd_sc_hd__nor2b_1
XFILLER_176_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7926_ fd._3223_ fd._3227_ fd._3229_ VGND VGND VPWR VPWR fd._3246_ sky130_fd_sc_hd__a21oi_1
XFILLER_108_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7857_ fd._3074_ fd._3038_ fd._3050_ fd._3060_ fd._1764_ VGND VGND VPWR VPWR fd._3170_
+ sky130_fd_sc_hd__a311o_1
XFILLER_195_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._6808_ fd._1842_ fd._1908_ VGND VGND VPWR VPWR fd._2016_ sky130_fd_sc_hd__nor2_1
Xfd._7788_ fd._2998_ fd._3008_ VGND VGND VPWR VPWR fd._3094_ sky130_fd_sc_hd__xnor2_1
XFILLER_254_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6739_ fd._1749_ fd._1939_ fd._1917_ VGND VGND VPWR VPWR fd._1940_ sky130_fd_sc_hd__mux2_1
XFILLER_208_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_259_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_1615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_283_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5070_ fd._3883_ fd._0103_ VGND VGND VPWR VPWR fd._0104_ sky130_fd_sc_hd__and2_1
XTAP_3573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5972_ fd._1092_ fd._1094_ fd._1095_ fd._1036_ VGND VGND VPWR VPWR fd._1096_ sky130_fd_sc_hd__nor4b_1
XFILLER_18_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4923_ fd._3675_ fd._3998_ VGND VGND VPWR VPWR fd._4017_ sky130_fd_sc_hd__or2_1
XFILLER_185_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7711_ fd._2998_ fd._3008_ fd._3006_ VGND VGND VPWR VPWR fd._3009_ sky130_fd_sc_hd__o21a_1
XFILLER_9_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._7642_ fd._2930_ fd._2932_ fd._2874_ VGND VGND VPWR VPWR fd._2933_ sky130_fd_sc_hd__mux2_1
Xfd._4854_ fd._3943_ fd._3784_ VGND VGND VPWR VPWR fd._3948_ sky130_fd_sc_hd__xnor2_1
XFILLER_220_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_project_wrapper_220 VGND VGND VPWR VPWR user_project_wrapper_220/HI la_data_out[98]
+ sky130_fd_sc_hd__conb_1
XFILLER_142_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_project_wrapper_231 VGND VGND VPWR VPWR user_project_wrapper_231/HI la_data_out[109]
+ sky130_fd_sc_hd__conb_1
XFILLER_114_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_242 VGND VGND VPWR VPWR user_project_wrapper_242/HI la_data_out[120]
+ sky130_fd_sc_hd__conb_1
XFILLER_154_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7573_ fd._2636_ fd._2658_ VGND VGND VPWR VPWR fd._2857_ sky130_fd_sc_hd__nand2_1
Xuser_project_wrapper_253 VGND VGND VPWR VPWR user_project_wrapper_253/HI wbs_ack_o
+ sky130_fd_sc_hd__conb_1
Xfd._4785_ fd._3626_ fd._3875_ fd._3878_ VGND VGND VPWR VPWR fd._3879_ sky130_fd_sc_hd__a21boi_2
Xuser_project_wrapper_264 VGND VGND VPWR VPWR user_project_wrapper_264/HI wbs_dat_o[10]
+ sky130_fd_sc_hd__conb_1
XFILLER_153_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_275 VGND VGND VPWR VPWR user_project_wrapper_275/HI wbs_dat_o[21]
+ sky130_fd_sc_hd__conb_1
Xfd._6524_ fd._0207_ fd._1699_ fd._1702_ VGND VGND VPWR VPWR fd._1703_ sky130_fd_sc_hd__mux2_2
XFILLER_114_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6455_ fd._1430_ fd._1503_ VGND VGND VPWR VPWR fd._1628_ sky130_fd_sc_hd__and2_1
XFILLER_155_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5406_ fd._0471_ fd._0473_ VGND VGND VPWR VPWR fd._0474_ sky130_fd_sc_hd__xnor2_1
XFILLER_116_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6386_ fd._1551_ fd._1403_ VGND VGND VPWR VPWR fd._1552_ sky130_fd_sc_hd__nor2_1
XFILLER_3_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_261_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8125_ fd.b\[25\] fd.a\[25\] VGND VGND VPWR VPWR fd._3440_ sky130_fd_sc_hd__and2b_1
XFILLER_228_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5337_ fd._0207_ fd._0200_ VGND VGND VPWR VPWR fd._0398_ sky130_fd_sc_hd__xnor2_1
XFILLER_243_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_247_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8056_ fd._3221_ fd._3230_ fd._3238_ fd._3235_ VGND VGND VPWR VPWR fd._3389_ sky130_fd_sc_hd__a31o_1
XFILLER_64_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5268_ fd._0319_ fd._0321_ VGND VGND VPWR VPWR fd._0322_ sky130_fd_sc_hd__xnor2_1
XFILLER_130_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7007_ fd._1632_ fd._2041_ fd._2234_ VGND VGND VPWR VPWR fd._2235_ sky130_fd_sc_hd__a21oi_1
Xfd._4219_ fd._0560_ fd._1473_ VGND VGND VPWR VPWR fd._1594_ sky130_fd_sc_hd__xnor2_1
XFILLER_247_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5199_ fd._4011_ fd._0129_ VGND VGND VPWR VPWR fd._0246_ sky130_fd_sc_hd__or2_1
XFILLER_212_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_1631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_9208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7909_ fd._1507_ fd._3226_ VGND VGND VPWR VPWR fd._3227_ sky130_fd_sc_hd__nand2_1
XFILLER_109_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_259_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout72 net73 VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__buf_2
XFILLER_50_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_276_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4570_ fd._3522_ fd._3541_ fd._3520_ VGND VGND VPWR VPWR fd._3664_ sky130_fd_sc_hd__o21a_1
XFILLER_237_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._6240_ fd._1349_ fd._1387_ fd._1388_ VGND VGND VPWR VPWR fd._1391_ sky130_fd_sc_hd__a21o_1
XFILLER_277_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_280_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6171_ fd._0786_ fd._1313_ VGND VGND VPWR VPWR fd._1315_ sky130_fd_sc_hd__nand2_1
XFILLER_225_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5122_ fd._0158_ fd._0159_ fd._0060_ fd._0160_ VGND VGND VPWR VPWR fd._0161_ sky130_fd_sc_hd__o31a_1
XTAP_4093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5053_ fd._4019_ fd._0084_ VGND VGND VPWR VPWR fd._0085_ sky130_fd_sc_hd__xnor2_1
XFILLER_233_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_261_1596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5955_ fd._1069_ fd._1076_ VGND VGND VPWR VPWR fd._1078_ sky130_fd_sc_hd__or2_1
XFILLER_179_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1670 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4906_ fd._3879_ fd._3954_ fd._3958_ VGND VGND VPWR VPWR fd._4000_ sky130_fd_sc_hd__nand3b_1
XFILLER_179_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._5886_ fd._0504_ fd._0999_ VGND VGND VPWR VPWR fd._1002_ sky130_fd_sc_hd__nand2_1
XFILLER_161_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4837_ fd._1352_ fd._3802_ VGND VGND VPWR VPWR fd._3931_ sky130_fd_sc_hd__and2_1
Xfd._7625_ fd._2780_ fd._2778_ VGND VGND VPWR VPWR fd._2915_ sky130_fd_sc_hd__nor2_1
XFILLER_115_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4768_ fd._3861_ VGND VGND VPWR VPWR fd._3862_ sky130_fd_sc_hd__inv_2
XFILLER_173_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7556_ fd._2836_ fd._2838_ VGND VGND VPWR VPWR fd._2839_ sky130_fd_sc_hd__and2_1
XFILLER_114_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6507_ fd._0967_ VGND VGND VPWR VPWR fd._1685_ sky130_fd_sc_hd__buf_6
XFILLER_134_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_275_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7487_ fd._1976_ VGND VGND VPWR VPWR fd._2763_ sky130_fd_sc_hd__buf_6
XFILLER_25_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4699_ fd._3791_ fd._3792_ VGND VGND VPWR VPWR fd._3793_ sky130_fd_sc_hd__or2_1
XFILLER_190_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_284_840 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6438_ fd._0343_ fd._1534_ VGND VGND VPWR VPWR fd._1609_ sky130_fd_sc_hd__nor2_1
XFILLER_25_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_283_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6369_ fd._1532_ VGND VGND VPWR VPWR fd._1533_ sky130_fd_sc_hd__buf_6
XFILLER_95_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8108_ fd._3424_ VGND VGND VPWR VPWR fd.mc\[21\] sky130_fd_sc_hd__buf_2
XFILLER_71_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_212_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8039_ fd._3096_ fd._3207_ VGND VGND VPWR VPWR fd._3370_ sky130_fd_sc_hd__nand2_1
XFILLER_266_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_252_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_9005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_8326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_277_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1590 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_259_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_1604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_236_ fd.c\[28\] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5740_ fd._0840_ VGND VGND VPWR VPWR fd._0841_ sky130_fd_sc_hd__inv_2
XFILLER_144_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_1610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5671_ fd._0601_ fd._0764_ fd._0672_ VGND VGND VPWR VPWR fd._0765_ sky130_fd_sc_hd__or3_1
XFILLER_143_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._4622_ fd.b\[11\] VGND VGND VPWR VPWR fd._3716_ sky130_fd_sc_hd__buf_6
Xfd._7410_ fd._2620_ fd._2670_ fd._2675_ VGND VGND VPWR VPWR fd._2678_ sky130_fd_sc_hd__and3_1
XFILLER_139_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7341_ fd._2411_ fd._2410_ VGND VGND VPWR VPWR fd._2602_ sky130_fd_sc_hd__nor2_1
Xfd._4553_ fd._0428_ fd._3502_ fd._3545_ VGND VGND VPWR VPWR fd._3647_ sky130_fd_sc_hd__a21o_1
XFILLER_170_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7272_ fd._2360_ VGND VGND VPWR VPWR fd._2526_ sky130_fd_sc_hd__inv_2
Xfd._4484_ fd._3565_ fd._3575_ fd._3577_ VGND VGND VPWR VPWR fd._3578_ sky130_fd_sc_hd__a21bo_1
XFILLER_152_1674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_272_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._6223_ fd._1195_ VGND VGND VPWR VPWR fd._1372_ sky130_fd_sc_hd__clkinv_2
XFILLER_37_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6154_ fd._1275_ fd._1237_ fd._1294_ VGND VGND VPWR VPWR fd._1296_ sky130_fd_sc_hd__and3_1
XFILLER_53_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5105_ fd._0141_ VGND VGND VPWR VPWR fd._0143_ sky130_fd_sc_hd__clkinv_4
XFILLER_111_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_263_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6085_ fd._1007_ fd._1032_ fd._1003_ VGND VGND VPWR VPWR fd._1221_ sky130_fd_sc_hd__o21ai_1
XFILLER_209_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5036_ fd._0060_ VGND VGND VPWR VPWR fd._0067_ sky130_fd_sc_hd__buf_6
XFILLER_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_267_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6987_ fd._2206_ fd._2211_ fd._1102_ VGND VGND VPWR VPWR fd._2213_ sky130_fd_sc_hd__a21o_1
XFILLER_105_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_257_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5938_ fd._1048_ fd._1052_ fd._1058_ VGND VGND VPWR VPWR fd._1059_ sky130_fd_sc_hd__o21bai_2
XFILLER_146_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5869_ fd._0981_ fd._0982_ VGND VGND VPWR VPWR fd._0983_ sky130_fd_sc_hd__nor2_1
XFILLER_162_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7608_ fd._2706_ fd._2895_ fd._2875_ VGND VGND VPWR VPWR fd._2896_ sky130_fd_sc_hd__mux2_1
XFILLER_161_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_255_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7539_ fd._2688_ fd._2810_ VGND VGND VPWR VPWR fd._2820_ sky130_fd_sc_hd__nor2_1
XFILLER_114_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_275_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_268_1547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_273_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_267_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_251_1584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_88 VGND VGND VPWR VPWR user_project_wrapper_88/HI io_oeb[10]
+ sky130_fd_sc_hd__conb_1
XFILLER_284_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_project_wrapper_99 VGND VGND VPWR VPWR user_project_wrapper_99/HI io_oeb[21]
+ sky130_fd_sc_hd__conb_1
XFILLER_216_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._6910_ fd._1986_ fd._2127_ VGND VGND VPWR VPWR fd._2128_ sky130_fd_sc_hd__xnor2_1
XFILLER_124_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7890_ fd._3205_ VGND VGND VPWR VPWR fd._3206_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_19_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6841_ fd._1846_ fd._2020_ fd._2051_ VGND VGND VPWR VPWR fd._2052_ sky130_fd_sc_hd__o21a_1
XFILLER_15_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_219_ fd.c\[11\] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
XFILLER_129_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6772_ fd._1397_ VGND VGND VPWR VPWR fd._1976_ sky130_fd_sc_hd__buf_6
XFILLER_128_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5723_ fd._0821_ fd._0636_ VGND VGND VPWR VPWR fd._0822_ sky130_fd_sc_hd__xnor2_1
XFILLER_183_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_256_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._5654_ fd._0653_ fd._0745_ VGND VGND VPWR VPWR fd._0746_ sky130_fd_sc_hd__nand2_1
XFILLER_143_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4605_ fd._3687_ fd._3694_ fd._3697_ fd._3698_ VGND VGND VPWR VPWR fd._3699_ sky130_fd_sc_hd__a31oi_4
XFILLER_217_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5585_ fd._0514_ fd._0521_ fd._0524_ VGND VGND VPWR VPWR fd._0671_ sky130_fd_sc_hd__and3_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_258_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_257_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._4536_ fd._2584_ fd._3568_ fd._3629_ VGND VGND VPWR VPWR fd._3630_ sky130_fd_sc_hd__o21ai_1
Xfd._7324_ fd._2326_ fd._2582_ VGND VGND VPWR VPWR fd._2583_ sky130_fd_sc_hd__xnor2_1
XFILLER_85_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_285_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_250_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7255_ fd._2324_ fd._2420_ fd._2506_ VGND VGND VPWR VPWR fd._2508_ sky130_fd_sc_hd__mux2_1
XFILLER_38_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4467_ fd._3439_ VGND VGND VPWR VPWR fd._3561_ sky130_fd_sc_hd__inv_2
XFILLER_239_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_272_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6206_ fd._1219_ fd._1224_ VGND VGND VPWR VPWR fd._1354_ sky130_fd_sc_hd__or2_1
XFILLER_39_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7186_ fd._2428_ fd._2431_ VGND VGND VPWR VPWR fd._2432_ sky130_fd_sc_hd__xnor2_1
XFILLER_54_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4398_ fd._0428_ fd._2111_ VGND VGND VPWR VPWR fd._3492_ sky130_fd_sc_hd__nor2_1
XFILLER_199_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_281_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6137_ fd._1118_ fd._1277_ VGND VGND VPWR VPWR fd._1278_ sky130_fd_sc_hd__nor2_1
XFILLER_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6068_ fd._1025_ fd._1201_ VGND VGND VPWR VPWR fd._1202_ sky130_fd_sc_hd__and2_1
XFILLER_0_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._5019_ fd._3957_ fd._0047_ VGND VGND VPWR VPWR fd._0048_ sky130_fd_sc_hd__nor2_1
XFILLER_221_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput38 net38 VGND VGND VPWR VPWR io_out[13] sky130_fd_sc_hd__buf_2
XFILLER_122_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput49 net49 VGND VGND VPWR VPWR io_out[23] sky130_fd_sc_hd__buf_2
XFILLER_270_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_276_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_281_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_279_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_253_1668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5370_ fd._0258_ fd._0433_ VGND VGND VPWR VPWR fd._0434_ sky130_fd_sc_hd__xnor2_1
XTAP_6573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4321_ fd._2694_ fd._2705_ VGND VGND VPWR VPWR fd._2716_ sky130_fd_sc_hd__or2b_1
XFILLER_255_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7040_ fd._2084_ fd._2088_ fd._2094_ VGND VGND VPWR VPWR fd._2271_ sky130_fd_sc_hd__o21a_1
XFILLER_75_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4252_ fd.b\[0\] fd.a\[0\] fd._1209_ VGND VGND VPWR VPWR fd._1957_ sky130_fd_sc_hd__and3_1
XFILLER_169_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4183_ fd.a\[22\] fd._4049_ VGND VGND VPWR VPWR fd._1198_ sky130_fd_sc_hd__and2_1
XFILLER_23_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_250_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_250_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7942_ fd._0768_ fd._3261_ VGND VGND VPWR VPWR fd._3263_ sky130_fd_sc_hd__nand2_1
XFILLER_15_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7873_ fd._3186_ VGND VGND VPWR VPWR fd._3187_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_129_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6824_ fd._2021_ fd._2026_ fd._2032_ VGND VGND VPWR VPWR fd._2033_ sky130_fd_sc_hd__a21o_1
XFILLER_15_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6755_ fd._1015_ VGND VGND VPWR VPWR fd._1958_ sky130_fd_sc_hd__buf_6
XFILLER_105_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5706_ fd._1341_ fd._0803_ VGND VGND VPWR VPWR fd._0804_ sky130_fd_sc_hd__and2_1
XFILLER_104_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6686_ fd._1878_ fd._1881_ VGND VGND VPWR VPWR fd._1882_ sky130_fd_sc_hd__nor2_1
XFILLER_158_1680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_258_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5637_ fd._0555_ fd._0727_ VGND VGND VPWR VPWR fd._0728_ sky130_fd_sc_hd__xnor2_1
XFILLER_131_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_258_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5568_ fd._0649_ fd._0650_ fd._0651_ VGND VGND VPWR VPWR fd._0652_ sky130_fd_sc_hd__mux2_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_1590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7307_ fd._2532_ fd._2538_ fd._2561_ fd._2563_ fd._2564_ VGND VGND VPWR VPWR fd._2565_
+ sky130_fd_sc_hd__a311o_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4519_ fd._3611_ fd._3612_ VGND VGND VPWR VPWR fd._3613_ sky130_fd_sc_hd__nand2_1
XFILLER_227_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5499_ fd._0573_ fd._0574_ fd._0452_ fd._0575_ VGND VGND VPWR VPWR fd._0576_ sky130_fd_sc_hd__a31o_1
XFILLER_6_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7238_ fd._2487_ fd._2488_ VGND VGND VPWR VPWR fd._2489_ sky130_fd_sc_hd__nor2_1
XFILLER_2_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_260_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_282_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7169_ fd._2126_ fd._2222_ VGND VGND VPWR VPWR fd._2413_ sky130_fd_sc_hd__nor2_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_257_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_268_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_274_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_1699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_1663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_264_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4870_ fd._3934_ fd._3803_ fd._3932_ VGND VGND VPWR VPWR fd._3964_ sky130_fd_sc_hd__nand3_1
XFILLER_201_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6540_ fd._1535_ fd._1612_ fd._1720_ VGND VGND VPWR VPWR fd._1721_ sky130_fd_sc_hd__mux2_1
XFILLER_113_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_1552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6471_ fd._4055_ VGND VGND VPWR VPWR fd._1645_ sky130_fd_sc_hd__buf_6
XFILLER_113_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._8210_ net74 net23 VGND VGND VPWR VPWR fd.a\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_256_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5422_ fd._3905_ fd._0490_ VGND VGND VPWR VPWR fd._0491_ sky130_fd_sc_hd__nor2_1
XTAP_7093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8141_ fd._3447_ fd._3455_ VGND VGND VPWR VPWR fd._3456_ sky130_fd_sc_hd__nor2_1
Xfd._5353_ fd._0214_ fd._0414_ fd._0270_ VGND VGND VPWR VPWR fd._0415_ sky130_fd_sc_hd__mux2_1
XFILLER_132_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4304_ fd._0714_ fd._2518_ VGND VGND VPWR VPWR fd._2529_ sky130_fd_sc_hd__xnor2_1
XTAP_5691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8072_ fd._2813_ fd._2877_ fd._3398_ VGND VGND VPWR VPWR fd._3402_ sky130_fd_sc_hd__mux2_2
XFILLER_76_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5284_ fd._3980_ fd._0300_ VGND VGND VPWR VPWR fd._0339_ sky130_fd_sc_hd__nand2_1
XFILLER_3_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_282_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_282_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4235_ fd._0318_ fd.a\[3\] VGND VGND VPWR VPWR fd._1770_ sky130_fd_sc_hd__nand2_1
XFILLER_235_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7023_ fd._2066_ fd._2103_ VGND VGND VPWR VPWR fd._2252_ sky130_fd_sc_hd__and2b_1
XFILLER_97_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_1657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_282_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4166_ fd._0164_ fd._0142_ VGND VGND VPWR VPWR fd._1011_ sky130_fd_sc_hd__or2b_1
XFILLER_251_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_264_1583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_264_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4097_ fd.b\[5\] VGND VGND VPWR VPWR fd._0252_ sky130_fd_sc_hd__buf_6
XFILLER_250_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7925_ fd._3220_ VGND VGND VPWR VPWR fd._3245_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_137_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7856_ fd._3075_ fd._3165_ fd._3168_ fd._2763_ VGND VGND VPWR VPWR fd._3169_ sky130_fd_sc_hd__a211o_1
XFILLER_34_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_258_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1554 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6807_ fd._2013_ fd._2014_ VGND VGND VPWR VPWR fd._2015_ sky130_fd_sc_hd__xnor2_1
XFILLER_129_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7787_ fd._1286_ fd._3092_ VGND VGND VPWR VPWR fd._3093_ sky130_fd_sc_hd__or2_1
Xfd._4999_ fd._3035_ VGND VGND VPWR VPWR fd._0026_ sky130_fd_sc_hd__buf_6
XFILLER_195_1655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_219_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_254_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6738_ fd._1937_ fd._1938_ VGND VGND VPWR VPWR fd._1939_ sky130_fd_sc_hd__xnor2_1
XFILLER_195_1688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_259_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6669_ fd._1859_ fd._1860_ fd._1861_ fd._1862_ VGND VGND VPWR VPWR fd._1863_ sky130_fd_sc_hd__o31a_1
XFILLER_132_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_1685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_273_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_274_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_230_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_272_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_269_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_277_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1690 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5971_ fd._1003_ fd._1007_ fd._1032_ fd._1037_ fd._1001_ VGND VGND VPWR VPWR fd._1095_
+ sky130_fd_sc_hd__o311a_1
XFILLER_119_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_28 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7710_ fd._3006_ fd._3007_ VGND VGND VPWR VPWR fd._3008_ sky130_fd_sc_hd__nand2_1
Xfd._4922_ fd._3883_ fd._3992_ VGND VGND VPWR VPWR fd._4016_ sky130_fd_sc_hd__or2_1
XFILLER_174_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7641_ fd._2931_ fd._2768_ VGND VGND VPWR VPWR fd._2932_ sky130_fd_sc_hd__xor2_1
XFILLER_127_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4853_ fd.b\[22\] VGND VGND VPWR VPWR fd._3947_ sky130_fd_sc_hd__buf_6
XFILLER_161_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_project_wrapper_210 VGND VGND VPWR VPWR user_project_wrapper_210/HI la_data_out[88]
+ sky130_fd_sc_hd__conb_1
Xuser_project_wrapper_221 VGND VGND VPWR VPWR user_project_wrapper_221/HI la_data_out[99]
+ sky130_fd_sc_hd__conb_1
XFILLER_182_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_project_wrapper_232 VGND VGND VPWR VPWR user_project_wrapper_232/HI la_data_out[110]
+ sky130_fd_sc_hd__conb_1
XFILLER_127_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_243 VGND VGND VPWR VPWR user_project_wrapper_243/HI la_data_out[121]
+ sky130_fd_sc_hd__conb_1
Xfd._7572_ fd._2853_ fd._2813_ fd._2854_ fd._2855_ VGND VGND VPWR VPWR fd._2856_ sky130_fd_sc_hd__a31o_1
XFILLER_5_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4784_ fd._3772_ fd._3783_ fd._3785_ fd._3877_ VGND VGND VPWR VPWR fd._3878_ sky130_fd_sc_hd__a31o_1
XFILLER_114_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_project_wrapper_254 VGND VGND VPWR VPWR user_project_wrapper_254/HI wbs_dat_o[0]
+ sky130_fd_sc_hd__conb_1
XFILLER_99_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_265 VGND VGND VPWR VPWR user_project_wrapper_265/HI wbs_dat_o[11]
+ sky130_fd_sc_hd__conb_1
Xuser_project_wrapper_276 VGND VGND VPWR VPWR user_project_wrapper_276/HI wbs_dat_o[22]
+ sky130_fd_sc_hd__conb_1
Xfd._6523_ fd._1700_ fd._1701_ VGND VGND VPWR VPWR fd._1702_ sky130_fd_sc_hd__xnor2_1
XFILLER_153_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_1382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6454_ fd._1618_ fd._1622_ fd._1625_ VGND VGND VPWR VPWR fd._1626_ sky130_fd_sc_hd__a21oi_4
XFILLER_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5405_ fd._0412_ fd._0401_ VGND VGND VPWR VPWR fd._0473_ sky130_fd_sc_hd__and2b_1
XFILLER_112_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6385_ fd._0312_ fd._1548_ VGND VGND VPWR VPWR fd._1551_ sky130_fd_sc_hd__nor2_1
XFILLER_151_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_256_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8124_ fd._3438_ VGND VGND VPWR VPWR fd.ec\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_55_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5336_ fd._0283_ fd._0387_ fd._0396_ VGND VGND VPWR VPWR fd._0397_ sky130_fd_sc_hd__a21o_1
XFILLER_7_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5267_ fd._0119_ fd._0320_ VGND VGND VPWR VPWR fd._0321_ sky130_fd_sc_hd__nor2_1
Xfd._8055_ fd._2863_ fd._3252_ VGND VGND VPWR VPWR fd._3388_ sky130_fd_sc_hd__nor2_1
XFILLER_247_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4218_ fd._1572_ VGND VGND VPWR VPWR fd._1583_ sky130_fd_sc_hd__inv_2
XFILLER_212_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7006_ fd._2233_ fd._2109_ VGND VGND VPWR VPWR fd._2234_ sky130_fd_sc_hd__and2_1
XFILLER_266_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5198_ fd._0125_ fd._0236_ VGND VGND VPWR VPWR fd._0245_ sky130_fd_sc_hd__nand2_1
XFILLER_169_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4149_ fd._0725_ fd._0747_ fd._0769_ fd._0813_ VGND VGND VPWR VPWR fd._0824_ sky130_fd_sc_hd__or4b_1
XFILLER_17_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7908_ fd._3042_ fd._3225_ fd._3077_ VGND VGND VPWR VPWR fd._3226_ sky130_fd_sc_hd__mux2_1
XFILLER_17_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7839_ fd._2944_ fd._2962_ VGND VGND VPWR VPWR fd._3150_ sky130_fd_sc_hd__xnor2_1
XTAP_8519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_273_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_258_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_273_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_259_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_246_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_274_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_251_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_280_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout73 net74 VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_4
XFILLER_204_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_276_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_269_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_1544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._6170_ fd._0786_ fd._1313_ VGND VGND VPWR VPWR fd._1314_ sky130_fd_sc_hd__or2_1
XFILLER_4_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5121_ fd._4032_ fd._0060_ VGND VGND VPWR VPWR fd._0160_ sky130_fd_sc_hd__nand2_1
XFILLER_225_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5052_ fd._4026_ fd._4024_ VGND VGND VPWR VPWR fd._0084_ sky130_fd_sc_hd__or2b_1
XFILLER_61_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5954_ fd._1088_ fd._1068_ VGND VGND VPWR VPWR fd._1076_ sky130_fd_sc_hd__nor2_1
XFILLER_105_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4905_ fd._3675_ fd._3998_ VGND VGND VPWR VPWR fd._3999_ sky130_fd_sc_hd__xnor2_1
XFILLER_220_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5885_ fd._0504_ fd._0999_ VGND VGND VPWR VPWR fd._1001_ sky130_fd_sc_hd__or2_1
XFILLER_122_1682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._7624_ fd._2776_ VGND VGND VPWR VPWR fd._2913_ sky130_fd_sc_hd__clkinv_2
XFILLER_255_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._4836_ fd._3813_ fd._3928_ fd._3929_ VGND VGND VPWR VPWR fd._3930_ sky130_fd_sc_hd__o21ba_1
XFILLER_192_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7555_ fd._2481_ fd._2835_ VGND VGND VPWR VPWR fd._2838_ sky130_fd_sc_hd__or2_1
Xfd._4767_ fd._0252_ fd._3860_ VGND VGND VPWR VPWR fd._3861_ sky130_fd_sc_hd__and2_1
XFILLER_170_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6506_ fd._1674_ fd._1681_ fd._1683_ VGND VGND VPWR VPWR fd._1684_ sky130_fd_sc_hd__o21bai_1
XFILLER_130_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7486_ fd._2670_ fd._2675_ fd._2761_ VGND VGND VPWR VPWR fd._2762_ sky130_fd_sc_hd__a21oi_1
Xfd._4698_ fd._3790_ fd._3751_ fd._3750_ fd._3633_ VGND VGND VPWR VPWR fd._3792_ sky130_fd_sc_hd__o211a_1
XFILLER_151_1322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6437_ fd._1543_ fd._1547_ fd._1599_ fd._1606_ fd._1607_ VGND VGND VPWR VPWR fd._1608_
+ sky130_fd_sc_hd__a41o_1
XFILLER_116_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_284_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6368_ fd._1513_ fd._1525_ fd._1531_ VGND VGND VPWR VPWR fd._1532_ sky130_fd_sc_hd__a21o_1
XFILLER_3_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8107_ fd._3626_ fd._3800_ fd._3189_ VGND VGND VPWR VPWR fd._3424_ sky130_fd_sc_hd__mux2_1
XFILLER_244_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._5319_ fd._0376_ fd._0377_ fd._0270_ VGND VGND VPWR VPWR fd._0378_ sky130_fd_sc_hd__mux2_1
XFILLER_243_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6299_ fd._1454_ fd._1455_ VGND VGND VPWR VPWR fd._1456_ sky130_fd_sc_hd__nor2_1
XFILLER_71_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._8038_ fd._2055_ fd._3368_ VGND VGND VPWR VPWR fd._3369_ sky130_fd_sc_hd__nand2_1
XFILLER_110_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_262_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_252_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_251_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_260_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_273_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_278_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_271_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_235_ fd.c\[27\] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_1
XFILLER_196_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5670_ fd._0482_ fd._0600_ VGND VGND VPWR VPWR fd._0764_ sky130_fd_sc_hd__and2_1
XTAP_8850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._4621_ fd._3655_ fd._3663_ fd._3710_ fd._3712_ fd._3714_ VGND VGND VPWR VPWR fd._3715_
+ sky130_fd_sc_hd__a311oi_2
XFILLER_139_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_8872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7340_ fd._2596_ fd._2599_ fd._2600_ VGND VGND VPWR VPWR fd._2601_ sky130_fd_sc_hd__a21oi_1
XFILLER_112_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4552_ fd.b\[14\] VGND VGND VPWR VPWR fd._3646_ sky130_fd_sc_hd__buf_6
XFILLER_65_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4483_ fd._1253_ fd._3571_ fd._3576_ VGND VGND VPWR VPWR fd._3577_ sky130_fd_sc_hd__a21o_1
XFILLER_152_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._7271_ fd._2367_ fd._2374_ fd._2383_ fd._2384_ VGND VGND VPWR VPWR fd._2525_ sky130_fd_sc_hd__a31o_1
XFILLER_46_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6222_ fd._1369_ fd._1370_ VGND VGND VPWR VPWR fd._1371_ sky130_fd_sc_hd__nor2_1
XFILLER_38_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6153_ fd._1237_ fd._1294_ fd._1275_ VGND VGND VPWR VPWR fd._1295_ sky130_fd_sc_hd__a21o_1
XFILLER_92_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5104_ fd._0090_ fd._0083_ VGND VGND VPWR VPWR fd._0141_ sky130_fd_sc_hd__or2b_1
XFILLER_209_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6084_ fd._0526_ VGND VGND VPWR VPWR fd._1219_ sky130_fd_sc_hd__buf_6
XFILLER_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5035_ fd._3972_ fd._0008_ fd._0063_ VGND VGND VPWR VPWR fd._0066_ sky130_fd_sc_hd__nand3_1
XFILLER_233_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6986_ fd._2206_ fd._2211_ VGND VGND VPWR VPWR fd._2212_ sky130_fd_sc_hd__or2_1
XFILLER_14_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5937_ fd._1053_ fd._1054_ fd._1057_ VGND VGND VPWR VPWR fd._1058_ sky130_fd_sc_hd__a21oi_1
XFILLER_107_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5868_ fd._0861_ fd._0863_ VGND VGND VPWR VPWR fd._0982_ sky130_fd_sc_hd__nand2_1
XFILLER_161_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7607_ fd._2894_ fd._2796_ VGND VGND VPWR VPWR fd._2895_ sky130_fd_sc_hd__xor2_1
XFILLER_115_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4819_ fd._3716_ fd._3912_ VGND VGND VPWR VPWR fd._3913_ sky130_fd_sc_hd__or2_1
XFILLER_216_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5799_ fd._0905_ fd._0686_ VGND VGND VPWR VPWR fd._0906_ sky130_fd_sc_hd__nor2_1
XFILLER_192_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7538_ fd._2684_ fd._2688_ fd._2810_ fd._2818_ fd._2680_ VGND VGND VPWR VPWR fd._2819_
+ sky130_fd_sc_hd__o311a_1
XTAP_5509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7469_ fd._2741_ VGND VGND VPWR VPWR fd._2743_ sky130_fd_sc_hd__inv_2
XTAP_4819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_262_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_273_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_1536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_251_1596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_263_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_262_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_78 VGND VGND VPWR VPWR user_project_wrapper_78/HI io_oeb[0]
+ sky130_fd_sc_hd__conb_1
XFILLER_28_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_89 VGND VGND VPWR VPWR user_project_wrapper_89/HI io_oeb[11]
+ sky130_fd_sc_hd__conb_1
XFILLER_147_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6840_ fd._2049_ fd._2050_ fd._1969_ VGND VGND VPWR VPWR fd._2051_ sky130_fd_sc_hd__or3_1
XFILLER_156_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_218_ fd.c\[10\] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6771_ fd._1969_ fd._1971_ fd._1974_ fd._1397_ VGND VGND VPWR VPWR fd._1975_ sky130_fd_sc_hd__a211o_1
XFILLER_237_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5722_ fd._0256_ VGND VGND VPWR VPWR fd._0821_ sky130_fd_sc_hd__buf_6
XFILLER_144_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_256_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5653_ fd._1275_ fd._0652_ VGND VGND VPWR VPWR fd._0745_ sky130_fd_sc_hd__nand2_1
XFILLER_28_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._4604_ fd.b\[3\] fd._3686_ VGND VGND VPWR VPWR fd._3698_ sky130_fd_sc_hd__nor2_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._5584_ fd._0668_ VGND VGND VPWR VPWR fd._0669_ sky130_fd_sc_hd__inv_2
XFILLER_174_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7323_ fd._2577_ fd._2579_ fd._2580_ fd._2581_ VGND VGND VPWR VPWR fd._2582_ sky130_fd_sc_hd__o31a_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4535_ fd._3565_ fd._3569_ VGND VGND VPWR VPWR fd._3629_ sky130_fd_sc_hd__nand2_1
XFILLER_257_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_250_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7254_ fd._2505_ VGND VGND VPWR VPWR fd._2506_ sky130_fd_sc_hd__buf_6
Xfd._4466_ fd._3422_ fd._3559_ VGND VGND VPWR VPWR fd._3560_ sky130_fd_sc_hd__nand2_1
XFILLER_26_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6205_ fd._1224_ VGND VGND VPWR VPWR fd._1353_ sky130_fd_sc_hd__clkinv_2
XFILLER_187_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_265_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7185_ fd._2429_ fd._2289_ VGND VGND VPWR VPWR fd._2431_ sky130_fd_sc_hd__nor2_1
XFILLER_93_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4397_ fd._1704_ fd._2078_ VGND VGND VPWR VPWR fd._3491_ sky130_fd_sc_hd__nor2_1
XFILLER_38_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6136_ fd._1249_ fd._1276_ fd._1246_ VGND VGND VPWR VPWR fd._1277_ sky130_fd_sc_hd__o21a_1
XFILLER_281_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6067_ fd._0638_ fd._1197_ VGND VGND VPWR VPWR fd._1201_ sky130_fd_sc_hd__nand2_1
XFILLER_185_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._5018_ fd._0044_ fd._3952_ fd._3950_ VGND VGND VPWR VPWR fd._0047_ sky130_fd_sc_hd__a21oi_1
XFILLER_210_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6969_ fd._2135_ fd._2139_ VGND VGND VPWR VPWR fd._2193_ sky130_fd_sc_hd__nand2_1
XFILLER_162_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput39 net39 VGND VGND VPWR VPWR io_out[14] sky130_fd_sc_hd__buf_2
XFILLER_192_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_276_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_257_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_260_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_260_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_281_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_234_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4320_ fd.b\[17\] fd._2683_ VGND VGND VPWR VPWR fd._2705_ sky130_fd_sc_hd__or2_1
XTAP_5862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4251_ fd.b\[0\] fd._1209_ fd.a\[0\] VGND VGND VPWR VPWR fd._1946_ sky130_fd_sc_hd__a21oi_1
XFILLER_208_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4182_ fd._0010_ fd._1132_ fd._1154_ fd._1176_ VGND VGND VPWR VPWR fd._1187_ sky130_fd_sc_hd__o31a_1
XFILLER_263_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_225_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_250_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._7941_ fd._1242_ fd._3242_ fd._3261_ fd._0768_ VGND VGND VPWR VPWR fd._3262_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_203_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7872_ fd._3184_ fd._3185_ VGND VGND VPWR VPWR fd._3186_ sky130_fd_sc_hd__nor2_1
XFILLER_15_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6823_ fd._2029_ fd._2031_ VGND VGND VPWR VPWR fd._2032_ sky130_fd_sc_hd__nor2_1
XFILLER_129_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6754_ fd._0450_ fd._1955_ VGND VGND VPWR VPWR fd._1956_ sky130_fd_sc_hd__nor2_1
XFILLER_144_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_264_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5705_ fd._0617_ fd._0647_ fd._0801_ VGND VGND VPWR VPWR fd._0803_ sky130_fd_sc_hd__mux2_1
Xfd._6685_ fd._1872_ fd._1877_ VGND VGND VPWR VPWR fd._1881_ sky130_fd_sc_hd__and2_1
XFILLER_144_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5636_ fd._0563_ fd._0561_ VGND VGND VPWR VPWR fd._0727_ sky130_fd_sc_hd__and2b_1
XFILLER_158_1692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_285_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5567_ fd._0614_ VGND VGND VPWR VPWR fd._0651_ sky130_fd_sc_hd__buf_6
XFILLER_274_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7306_ fd._2141_ fd._2530_ VGND VGND VPWR VPWR fd._2564_ sky130_fd_sc_hd__and2_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4518_ fd.b\[22\] fd._3610_ VGND VGND VPWR VPWR fd._3612_ sky130_fd_sc_hd__nand2_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5498_ fd._0372_ fd._0452_ VGND VGND VPWR VPWR fd._0575_ sky130_fd_sc_hd__nor2_1
XFILLER_227_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7237_ fd._2481_ fd._2486_ VGND VGND VPWR VPWR fd._2488_ sky130_fd_sc_hd__nor2_1
XFILLER_22_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4449_ fd._3522_ fd._3541_ fd._3542_ fd._3520_ VGND VGND VPWR VPWR fd._3543_ sky130_fd_sc_hd__o211a_1
XFILLER_54_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7168_ fd._2404_ fd._2410_ fd._2411_ VGND VGND VPWR VPWR fd._2412_ sky130_fd_sc_hd__o21bai_1
XFILLER_54_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6119_ fd._1256_ fd._1257_ VGND VGND VPWR VPWR fd._1258_ sky130_fd_sc_hd__nand2_1
XFILLER_263_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7099_ fd._2140_ fd._2195_ fd._2134_ VGND VGND VPWR VPWR fd._2336_ sky130_fd_sc_hd__o21a_1
XFILLER_41_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_1614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_276_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_260_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._6470_ fd._1631_ fd._1637_ fd._1642_ fd._1643_ VGND VGND VPWR VPWR fd._1644_ sky130_fd_sc_hd__a211o_2
XFILLER_218_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5421_ fd._0488_ VGND VGND VPWR VPWR fd._0490_ sky130_fd_sc_hd__inv_2
XTAP_7083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_268_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8140_ fd._3453_ fd._3454_ VGND VGND VPWR VPWR fd._3455_ sky130_fd_sc_hd__nor2_1
XTAP_6382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5352_ fd._0272_ fd._0218_ VGND VGND VPWR VPWR fd._0414_ sky130_fd_sc_hd__xnor2_1
XTAP_6393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_255_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4303_ fd._0769_ fd._2430_ fd._0747_ VGND VGND VPWR VPWR fd._2518_ sky130_fd_sc_hd__o21bai_1
XFILLER_208_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._8071_ fd._3401_ VGND VGND VPWR VPWR fd.mc\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_97_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5283_ fd._3658_ fd._0335_ VGND VGND VPWR VPWR fd._0338_ sky130_fd_sc_hd__nor2_1
XFILLER_212_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_270_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7022_ fd._2075_ fd._2102_ fd._2073_ VGND VGND VPWR VPWR fd._2251_ sky130_fd_sc_hd__o21a_1
XTAP_4991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4234_ fd._0252_ fd._1748_ VGND VGND VPWR VPWR fd._1759_ sky130_fd_sc_hd__nand2_1
XFILLER_224_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_250_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4165_ fd._0989_ VGND VGND VPWR VPWR fd._1000_ sky130_fd_sc_hd__clkinv_4
XFILLER_51_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_259_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_260_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._4096_ fd.a\[5\] fd.b\[5\] VGND VGND VPWR VPWR fd._0241_ sky130_fd_sc_hd__nor2b_1
XFILLER_143_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7924_ fd._1242_ fd._3242_ VGND VGND VPWR VPWR fd._3243_ sky130_fd_sc_hd__or2_1
XFILLER_52_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_223_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7855_ fd._3021_ fd._3039_ fd._3051_ fd._3061_ fd._3166_ VGND VGND VPWR VPWR fd._3168_
+ sky130_fd_sc_hd__o311a_1
XFILLER_176_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6806_ fd._1661_ fd._1918_ VGND VGND VPWR VPWR fd._2014_ sky130_fd_sc_hd__xnor2_1
XFILLER_121_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_1634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7786_ fd._3014_ fd._3091_ fd._3077_ VGND VGND VPWR VPWR fd._3092_ sky130_fd_sc_hd__mux2_1
XFILLER_69_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4998_ fd._0016_ fd._0023_ fd._0024_ VGND VGND VPWR VPWR fd._0025_ sky130_fd_sc_hd__a21oi_1
XFILLER_145_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6737_ fd._1750_ fd._1775_ VGND VGND VPWR VPWR fd._1938_ sky130_fd_sc_hd__and2b_1
XFILLER_160_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._6668_ fd._1664_ fd._1861_ VGND VGND VPWR VPWR fd._1862_ sky130_fd_sc_hd__nand2_1
XFILLER_144_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_258_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5619_ fd._0700_ fd._0706_ fd._0707_ VGND VGND VPWR VPWR fd._0708_ sky130_fd_sc_hd__o21ba_1
XFILLER_86_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1588 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6599_ fd._1785_ VGND VGND VPWR VPWR fd._1786_ sky130_fd_sc_hd__inv_2
XFILLER_100_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_274_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8269_ net68 net22 VGND VGND VPWR VPWR fd.b\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5970_ fd._1089_ fd._1093_ VGND VGND VPWR VPWR fd._1094_ sky130_fd_sc_hd__nand2_1
XFILLER_13_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._4921_ fd._4005_ fd._4010_ fd._4013_ fd._4014_ VGND VGND VPWR VPWR fd._4015_ sky130_fd_sc_hd__o31a_1
XFILLER_201_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7640_ fd._2769_ fd._2750_ VGND VGND VPWR VPWR fd._2931_ sky130_fd_sc_hd__or2b_1
Xfd._4852_ fd._3766_ fd._3945_ fd._3800_ VGND VGND VPWR VPWR fd._3946_ sky130_fd_sc_hd__mux2_1
Xuser_project_wrapper_200 VGND VGND VPWR VPWR user_project_wrapper_200/HI la_data_out[78]
+ sky130_fd_sc_hd__conb_1
XFILLER_86_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_211 VGND VGND VPWR VPWR user_project_wrapper_211/HI la_data_out[89]
+ sky130_fd_sc_hd__conb_1
XFILLER_160_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_222 VGND VGND VPWR VPWR user_project_wrapper_222/HI la_data_out[100]
+ sky130_fd_sc_hd__conb_1
XFILLER_142_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7571_ fd._2667_ fd._2813_ VGND VGND VPWR VPWR fd._2855_ sky130_fd_sc_hd__nor2_1
Xuser_project_wrapper_233 VGND VGND VPWR VPWR user_project_wrapper_233/HI la_data_out[111]
+ sky130_fd_sc_hd__conb_1
Xfd._4783_ fd._3695_ fd._3876_ fd._3696_ VGND VGND VPWR VPWR fd._3877_ sky130_fd_sc_hd__o21ai_1
XFILLER_182_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_project_wrapper_244 VGND VGND VPWR VPWR user_project_wrapper_244/HI la_data_out[122]
+ sky130_fd_sc_hd__conb_1
XFILLER_153_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_project_wrapper_255 VGND VGND VPWR VPWR user_project_wrapper_255/HI wbs_dat_o[1]
+ sky130_fd_sc_hd__conb_1
Xuser_project_wrapper_266 VGND VGND VPWR VPWR user_project_wrapper_266/HI wbs_dat_o[12]
+ sky130_fd_sc_hd__conb_1
Xfd._6522_ fd._1431_ fd._1438_ VGND VGND VPWR VPWR fd._1701_ sky130_fd_sc_hd__xnor2_1
XFILLER_4_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_277 VGND VGND VPWR VPWR user_project_wrapper_277/HI wbs_dat_o[23]
+ sky130_fd_sc_hd__conb_1
XFILLER_218_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_1359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6453_ fd._1623_ fd._1624_ fd._1520_ VGND VGND VPWR VPWR fd._1625_ sky130_fd_sc_hd__mux2_1
XFILLER_68_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5404_ fd._0394_ fd._0470_ fd._0393_ VGND VGND VPWR VPWR fd._0471_ sky130_fd_sc_hd__a21bo_1
XFILLER_190_1586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_261_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6384_ fd._1383_ fd._1390_ fd._1401_ fd._1402_ VGND VGND VPWR VPWR fd._1549_ sky130_fd_sc_hd__a31o_1
XTAP_6190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8123_ fd._3436_ fd._3437_ VGND VGND VPWR VPWR fd._3438_ sky130_fd_sc_hd__or2_1
XFILLER_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_256_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5335_ fd._0393_ fd._0394_ VGND VGND VPWR VPWR fd._0396_ sky130_fd_sc_hd__nand2_1
XFILLER_209_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_255_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8054_ fd._3385_ fd._3381_ fd._3375_ VGND VGND VPWR VPWR fd._3386_ sky130_fd_sc_hd__a21bo_1
XFILLER_97_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5266_ fd._3869_ fd._0118_ VGND VGND VPWR VPWR fd._0320_ sky130_fd_sc_hd__nor2_1
XFILLER_3_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_247_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7005_ fd._2063_ fd._2108_ VGND VGND VPWR VPWR fd._2233_ sky130_fd_sc_hd__or2_1
Xfd._4217_ fd.b\[11\] fd._1561_ VGND VGND VPWR VPWR fd._1572_ sky130_fd_sc_hd__nand2_1
XFILLER_251_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5197_ fd._0227_ fd._0243_ fd._0234_ fd._0062_ VGND VGND VPWR VPWR fd._0244_ sky130_fd_sc_hd__o211ai_4
XFILLER_149_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4148_ fd._0791_ fd._0802_ VGND VGND VPWR VPWR fd._0813_ sky130_fd_sc_hd__and2b_1
XFILLER_71_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4079_ fd.b\[16\] fd._0043_ VGND VGND VPWR VPWR fd._0054_ sky130_fd_sc_hd__nor2_1
XFILLER_260_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7907_ fd._3217_ fd._3224_ VGND VGND VPWR VPWR fd._3225_ sky130_fd_sc_hd__or2_1
XFILLER_137_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7838_ fd._3147_ fd._3148_ VGND VGND VPWR VPWR fd._3149_ sky130_fd_sc_hd__nand2_1
XFILLER_121_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_258_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_273_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7769_ fd._2887_ fd._2893_ fd._3018_ fd._2885_ VGND VGND VPWR VPWR fd._3073_ sky130_fd_sc_hd__o31a_1
XFILLER_258_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_279_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_1328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_254_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_259_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_261_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_251_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_265_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_261_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout74 net75 VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_4
XFILLER_156_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_276_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_272_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_276_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_269_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_1583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_250_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_1556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5120_ fd._3982_ fd._4028_ fd._0157_ VGND VGND VPWR VPWR fd._0159_ sky130_fd_sc_hd__a21oi_1
XTAP_4073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_283_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5051_ fd._3469_ fd._0082_ VGND VGND VPWR VPWR fd._0083_ sky130_fd_sc_hd__or2_1
XFILLER_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_283_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5953_ fd._0479_ fd._1061_ VGND VGND VPWR VPWR fd._1075_ sky130_fd_sc_hd__and2_1
XFILLER_174_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4904_ fd._3873_ fd._3997_ fd._3959_ VGND VGND VPWR VPWR fd._3998_ sky130_fd_sc_hd__mux2_1
XFILLER_174_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5884_ fd._0809_ fd._0994_ fd._0998_ VGND VGND VPWR VPWR fd._0999_ sky130_fd_sc_hd__mux2_1
XFILLER_220_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_1694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7623_ fd._2566_ fd._2911_ VGND VGND VPWR VPWR fd._2912_ sky130_fd_sc_hd__or2_1
Xfd._4835_ fd._3580_ fd._3807_ VGND VGND VPWR VPWR fd._3929_ sky130_fd_sc_hd__nor2_1
XFILLER_127_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7554_ fd._2481_ fd._2835_ VGND VGND VPWR VPWR fd._2836_ sky130_fd_sc_hd__nand2_1
Xfd._4766_ fd._3859_ fd._3679_ fd._3787_ VGND VGND VPWR VPWR fd._3860_ sky130_fd_sc_hd__mux2_1
XFILLER_114_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_272_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._6505_ fd._1319_ fd._1680_ VGND VGND VPWR VPWR fd._1683_ sky130_fd_sc_hd__and2_1
XFILLER_272_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7485_ fd._1211_ fd._2753_ VGND VGND VPWR VPWR fd._2761_ sky130_fd_sc_hd__xnor2_1
XFILLER_114_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4697_ fd._3633_ fd._3750_ fd._3751_ fd._3790_ VGND VGND VPWR VPWR fd._3791_ sky130_fd_sc_hd__a211oi_1
XFILLER_130_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6436_ fd._1604_ fd._1541_ fd._1603_ VGND VGND VPWR VPWR fd._1607_ sky130_fd_sc_hd__a21oi_1
XFILLER_151_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6367_ fd._1520_ fd._1522_ fd._1530_ VGND VGND VPWR VPWR fd._1531_ sky130_fd_sc_hd__o21ai_1
XFILLER_95_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8106_ fd._3423_ VGND VGND VPWR VPWR fd.mc\[20\] sky130_fd_sc_hd__buf_2
XFILLER_243_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5318_ fd._0181_ fd._0177_ VGND VGND VPWR VPWR fd._0377_ sky130_fd_sc_hd__xnor2_1
XFILLER_37_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6298_ fd._0343_ fd._1453_ VGND VGND VPWR VPWR fd._1455_ sky130_fd_sc_hd__and2_1
XFILLER_243_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8037_ fd._3098_ fd._3367_ fd._3240_ VGND VGND VPWR VPWR fd._3368_ sky130_fd_sc_hd__mux2_1
XFILLER_52_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5249_ fd._3980_ fd._0300_ VGND VGND VPWR VPWR fd._0301_ sky130_fd_sc_hd__or2_1
XFILLER_24_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_267_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_262_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_264_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_1527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_234_ fd.c\[26\] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_1
XFILLER_156_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4620_ fd._3713_ VGND VGND VPWR VPWR fd._3714_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_276_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._4551_ fd._2584_ fd._3644_ VGND VGND VPWR VPWR fd._3645_ sky130_fd_sc_hd__or2_1
XFILLER_151_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7270_ fd._2359_ VGND VGND VPWR VPWR fd._2524_ sky130_fd_sc_hd__clkinv_2
Xfd._4482_ fd._2584_ fd._3568_ fd._3571_ fd._1253_ VGND VGND VPWR VPWR fd._3576_ sky130_fd_sc_hd__o22a_1
XFILLER_113_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6221_ fd._1178_ fd._1368_ VGND VGND VPWR VPWR fd._1370_ sky130_fd_sc_hd__nor2_1
XFILLER_66_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6152_ fd._1241_ fd._1283_ fd._1289_ fd._1292_ fd._1293_ VGND VGND VPWR VPWR fd._1294_
+ sky130_fd_sc_hd__a311o_1
XFILLER_4_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_280_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5103_ fd._3708_ fd._0139_ VGND VGND VPWR VPWR fd._0140_ sky130_fd_sc_hd__nor2_1
XFILLER_34_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6083_ fd._1185_ fd._1189_ fd._1216_ fd._1217_ VGND VGND VPWR VPWR fd._1218_ sky130_fd_sc_hd__a31o_1
XTAP_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_1638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5034_ fd._3972_ fd._0008_ fd._0063_ VGND VGND VPWR VPWR fd._0064_ sky130_fd_sc_hd__a21o_1
XFILLER_244_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_267_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6985_ fd._1923_ fd._2209_ fd._2116_ VGND VGND VPWR VPWR fd._2211_ sky130_fd_sc_hd__mux2_1
XFILLER_179_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5936_ fd._0850_ fd._1056_ VGND VGND VPWR VPWR fd._1057_ sky130_fd_sc_hd__xnor2_1
XFILLER_88_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5867_ fd._0869_ fd._0980_ VGND VGND VPWR VPWR fd._0981_ sky130_fd_sc_hd__nand2_1
XFILLER_146_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_1688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4818_ fd._3911_ fd._3650_ fd._3787_ VGND VGND VPWR VPWR fd._3912_ sky130_fd_sc_hd__mux2_1
Xfd._7606_ fd._2713_ fd._2794_ fd._2797_ VGND VGND VPWR VPWR fd._2894_ sky130_fd_sc_hd__o21ai_1
XFILLER_157_1554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5798_ fd._0526_ fd._0675_ VGND VGND VPWR VPWR fd._0905_ sky130_fd_sc_hd__and2_1
XFILLER_115_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_283_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_255_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7537_ fd._2816_ fd._2817_ VGND VGND VPWR VPWR fd._2818_ sky130_fd_sc_hd__nor2_1
XFILLER_130_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4749_ fd._3707_ fd._3842_ VGND VGND VPWR VPWR fd._3843_ sky130_fd_sc_hd__nand2_1
XFILLER_170_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7468_ fd._2533_ fd._2741_ VGND VGND VPWR VPWR fd._2742_ sky130_fd_sc_hd__nand2_1
XTAP_4809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_275_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_257_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6419_ fd._1584_ fd._1587_ fd._1532_ VGND VGND VPWR VPWR fd._1588_ sky130_fd_sc_hd__mux2_1
XFILLER_99_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7399_ fd._2660_ fd._2495_ VGND VGND VPWR VPWR fd._2666_ sky130_fd_sc_hd__xnor2_1
XFILLER_257_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_283_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_281_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_8103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_8147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_267_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_project_wrapper_79 VGND VGND VPWR VPWR user_project_wrapper_79/HI io_oeb[1]
+ sky130_fd_sc_hd__conb_1
XFILLER_28_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_217_ fd.c\[9\] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_1
Xfd._6770_ fd._1821_ fd._1835_ fd._1915_ fd._1973_ VGND VGND VPWR VPWR fd._1974_ sky130_fd_sc_hd__a31oi_1
XFILLER_15_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5721_ fd._0632_ fd._0631_ VGND VGND VPWR VPWR fd._0820_ sky130_fd_sc_hd__or2_1
XFILLER_156_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5652_ fd._0739_ fd._0743_ VGND VGND VPWR VPWR fd._0744_ sky130_fd_sc_hd__xnor2_1
XTAP_8670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._4603_ fd.b\[2\] fd._3693_ fd._3696_ VGND VGND VPWR VPWR fd._3697_ sky130_fd_sc_hd__o21ai_2
XFILLER_112_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._5583_ fd._0666_ fd._0667_ VGND VGND VPWR VPWR fd._0668_ sky130_fd_sc_hd__or2_1
XFILLER_152_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7322_ fd._2338_ fd._2577_ VGND VGND VPWR VPWR fd._2581_ sky130_fd_sc_hd__nand2_1
XFILLER_112_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4534_ fd._1352_ fd._3627_ VGND VGND VPWR VPWR fd._3628_ sky130_fd_sc_hd__or2_1
XTAP_7991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_273_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7253_ fd._2498_ fd._2504_ VGND VGND VPWR VPWR fd._2505_ sky130_fd_sc_hd__nand2_4
XFILLER_38_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4465_ fd.b\[12\] fd._3416_ VGND VGND VPWR VPWR fd._3559_ sky130_fd_sc_hd__nand2_1
XFILLER_250_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6204_ fd._1350_ VGND VGND VPWR VPWR fd._1351_ sky130_fd_sc_hd__clkinv_2
XFILLER_113_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7184_ fd._1286_ fd._2260_ VGND VGND VPWR VPWR fd._2429_ sky130_fd_sc_hd__and2_1
XFILLER_54_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_265_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4396_ fd._3469_ fd._3489_ VGND VGND VPWR VPWR fd._3490_ sky130_fd_sc_hd__or2_1
XFILLER_281_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6135_ fd._1267_ fd._1273_ fd._1274_ VGND VGND VPWR VPWR fd._1276_ sky130_fd_sc_hd__a21oi_1
XFILLER_187_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_281_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6066_ fd._0632_ fd._1027_ VGND VGND VPWR VPWR fd._1200_ sky130_fd_sc_hd__or2_1
XFILLER_62_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_263_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._5017_ fd._3949_ fd._0045_ fd._3961_ VGND VGND VPWR VPWR fd._0046_ sky130_fd_sc_hd__mux2_1
XFILLER_90_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6968_ fd._2165_ fd._2174_ fd._2189_ fd._2190_ fd._2191_ VGND VGND VPWR VPWR fd._2192_
+ sky130_fd_sc_hd__o311a_1
XFILLER_124_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5919_ fd._1036_ fd._1037_ VGND VGND VPWR VPWR fd._1038_ sky130_fd_sc_hd__nand2_1
XFILLER_200_1463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6899_ fd._2115_ VGND VGND VPWR VPWR fd._2116_ sky130_fd_sc_hd__buf_6
XFILLER_227_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_281_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_255_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4250_ fd.b\[2\] fd._1924_ VGND VGND VPWR VPWR fd._1935_ sky130_fd_sc_hd__nand2_1
XTAP_5896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._4181_ fd._1165_ fd.a\[21\] VGND VGND VPWR VPWR fd._1176_ sky130_fd_sc_hd__or2_1
XFILLER_78_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7940_ fd._3078_ fd._3260_ fd._3241_ VGND VGND VPWR VPWR fd._3261_ sky130_fd_sc_hd__mux2_1
XFILLER_30_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7871_ fd._2566_ fd._3183_ VGND VGND VPWR VPWR fd._3185_ sky130_fd_sc_hd__nor2_1
XFILLER_15_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6822_ fd._1830_ fd._2027_ fd._1969_ fd._2030_ VGND VGND VPWR VPWR fd._2031_ sky130_fd_sc_hd__o211a_1
XFILLER_30_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6753_ fd._1950_ fd._1954_ fd._1917_ VGND VGND VPWR VPWR fd._1955_ sky130_fd_sc_hd__mux2_1
XFILLER_183_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5704_ fd._0781_ fd._0794_ fd._0796_ fd._0800_ VGND VGND VPWR VPWR fd._0801_ sky130_fd_sc_hd__a211o_4
XFILLER_176_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6684_ fd._1878_ VGND VGND VPWR VPWR fd._1879_ sky130_fd_sc_hd__inv_2
XTAP_9190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5635_ fd._3646_ VGND VGND VPWR VPWR fd._0726_ sky130_fd_sc_hd__buf_6
XFILLER_113_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5566_ fd._0579_ fd._0584_ VGND VGND VPWR VPWR fd._0650_ sky130_fd_sc_hd__xor2_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4517_ fd.b\[22\] fd._3610_ VGND VGND VPWR VPWR fd._3611_ sky130_fd_sc_hd__or2_1
XFILLER_189_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7305_ fd._1219_ fd._2522_ VGND VGND VPWR VPWR fd._2563_ sky130_fd_sc_hd__nor2_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5497_ fd._0369_ fd._0374_ VGND VGND VPWR VPWR fd._0574_ sky130_fd_sc_hd__or2_1
XFILLER_117_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7236_ fd._2481_ fd._2486_ VGND VGND VPWR VPWR fd._2487_ sky130_fd_sc_hd__and2_1
XFILLER_94_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4448_ fd._0252_ fd._3512_ VGND VGND VPWR VPWR fd._3542_ sky130_fd_sc_hd__or2_1
XFILLER_187_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7167_ fd._1661_ fd._2409_ VGND VGND VPWR VPWR fd._2411_ sky130_fd_sc_hd__and2_1
Xfd._4379_ fd._2375_ fd._3343_ fd._3211_ VGND VGND VPWR VPWR fd._3354_ sky130_fd_sc_hd__a21bo_1
XFILLER_226_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6118_ fd._1102_ fd._1255_ VGND VGND VPWR VPWR fd._1257_ sky130_fd_sc_hd__or2_1
XFILLER_39_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_267_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._7098_ fd._2333_ fd._2334_ VGND VGND VPWR VPWR fd._2335_ sky130_fd_sc_hd__nand2_1
XFILLER_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6049_ fd._1007_ fd._1031_ VGND VGND VPWR VPWR fd._1181_ sky130_fd_sc_hd__nor2_1
XFILLER_165_1675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_263_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_281_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_1704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_268_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5420_ fd._0343_ fd._0488_ VGND VGND VPWR VPWR fd._0489_ sky130_fd_sc_hd__nor2_1
XFILLER_214_1407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5351_ fd._0397_ fd._0402_ fd._0411_ fd._0412_ VGND VGND VPWR VPWR fd._0413_ sky130_fd_sc_hd__a211oi_2
XTAP_6383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_255_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4302_ fd.a\[14\] VGND VGND VPWR VPWR fd._2507_ sky130_fd_sc_hd__clkinv_2
XTAP_5671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._8070_ fd._2877_ fd._3077_ fd._3398_ VGND VGND VPWR VPWR fd._3401_ sky130_fd_sc_hd__mux2_1
XFILLER_76_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5282_ fd._0089_ fd._0295_ VGND VGND VPWR VPWR fd._0337_ sky130_fd_sc_hd__xnor2_1
XTAP_5693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_264_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._7021_ fd._2239_ fd._2245_ fd._2249_ VGND VGND VPWR VPWR fd._2250_ sky130_fd_sc_hd__a21oi_4
XTAP_4970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4233_ fd._1715_ fd._1737_ fd._1209_ VGND VGND VPWR VPWR fd._1748_ sky130_fd_sc_hd__mux2_1
XFILLER_209_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._4164_ fd._0054_ fd._0978_ VGND VGND VPWR VPWR fd._0989_ sky130_fd_sc_hd__nor2_1
XFILLER_264_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_250_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_259_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4095_ fd._0219_ fd.a\[4\] VGND VGND VPWR VPWR fd._0230_ sky130_fd_sc_hd__xnor2_1
XFILLER_250_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7923_ fd._3065_ fd._3215_ fd._3241_ VGND VGND VPWR VPWR fd._3242_ sky130_fd_sc_hd__mux2_1
XFILLER_143_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7854_ fd._1970_ fd._2877_ VGND VGND VPWR VPWR fd._3166_ sky130_fd_sc_hd__nand2_1
XFILLER_125_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6805_ fd._2005_ fd._2010_ fd._2011_ VGND VGND VPWR VPWR fd._2013_ sky130_fd_sc_hd__a21oi_1
XFILLER_145_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4997_ fd._1352_ fd._0022_ VGND VGND VPWR VPWR fd._0024_ sky130_fd_sc_hd__and2_1
XFILLER_144_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7785_ fd._3009_ fd._3089_ VGND VGND VPWR VPWR fd._3091_ sky130_fd_sc_hd__xnor2_1
XFILLER_69_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6736_ fd._1934_ fd._1936_ fd._1774_ VGND VGND VPWR VPWR fd._1937_ sky130_fd_sc_hd__a21bo_1
XFILLER_208_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_271_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6667_ fd._1626_ fd._1644_ fd._1718_ VGND VGND VPWR VPWR fd._1861_ sky130_fd_sc_hd__and3_1
XFILLER_99_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_1676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_271_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5618_ fd._3905_ fd._0705_ VGND VGND VPWR VPWR fd._0707_ sky130_fd_sc_hd__and2_1
XFILLER_8_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6598_ fd._1783_ fd._1784_ VGND VGND VPWR VPWR fd._1785_ sky130_fd_sc_hd__nor2_1
XFILLER_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5549_ fd._0437_ fd._0465_ fd._0481_ fd._0612_ VGND VGND VPWR VPWR fd._0631_ sky130_fd_sc_hd__and4_1
XFILLER_150_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_255_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8268_ net68 net21 VGND VGND VPWR VPWR fd.b\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_227_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7219_ fd._2297_ fd._2303_ fd._2302_ VGND VGND VPWR VPWR fd._2468_ sky130_fd_sc_hd__o21bai_1
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8199_ net66 fd.ec\[0\] VGND VGND VPWR VPWR fd.c\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_269_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_276_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_265_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_250_1629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_260_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4920_ fd._4000_ fd._4004_ fd._3869_ VGND VGND VPWR VPWR fd._4014_ sky130_fd_sc_hd__a21o_1
XFILLER_174_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._4851_ fd._3781_ fd._3944_ VGND VGND VPWR VPWR fd._3945_ sky130_fd_sc_hd__xnor2_1
XFILLER_127_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_project_wrapper_201 VGND VGND VPWR VPWR user_project_wrapper_201/HI la_data_out[79]
+ sky130_fd_sc_hd__conb_1
XFILLER_182_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_212 VGND VGND VPWR VPWR user_project_wrapper_212/HI la_data_out[90]
+ sky130_fd_sc_hd__conb_1
XFILLER_255_1507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_223 VGND VGND VPWR VPWR user_project_wrapper_223/HI la_data_out[101]
+ sky130_fd_sc_hd__conb_1
Xfd._4782_ fd._3537_ fd._3626_ VGND VGND VPWR VPWR fd._3876_ sky130_fd_sc_hd__or2_1
Xfd._7570_ fd._2852_ fd._2668_ VGND VGND VPWR VPWR fd._2854_ sky130_fd_sc_hd__or2_1
Xuser_project_wrapper_234 VGND VGND VPWR VPWR user_project_wrapper_234/HI la_data_out[112]
+ sky130_fd_sc_hd__conb_1
XFILLER_126_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_245 VGND VGND VPWR VPWR user_project_wrapper_245/HI la_data_out[123]
+ sky130_fd_sc_hd__conb_1
XFILLER_5_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_project_wrapper_256 VGND VGND VPWR VPWR user_project_wrapper_256/HI wbs_dat_o[2]
+ sky130_fd_sc_hd__conb_1
Xfd._6521_ fd._1499_ fd._1496_ fd._1617_ VGND VGND VPWR VPWR fd._1700_ sky130_fd_sc_hd__nand3b_1
XFILLER_175_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_267 VGND VGND VPWR VPWR user_project_wrapper_267/HI wbs_dat_o[13]
+ sky130_fd_sc_hd__conb_1
Xuser_project_wrapper_278 VGND VGND VPWR VPWR user_project_wrapper_278/HI wbs_dat_o[24]
+ sky130_fd_sc_hd__conb_1
XFILLER_142_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_268_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6452_ fd._1530_ fd._1623_ VGND VGND VPWR VPWR fd._1624_ sky130_fd_sc_hd__nor2_1
XFILLER_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5403_ fd._0283_ fd._0387_ VGND VGND VPWR VPWR fd._0470_ sky130_fd_sc_hd__nand2_1
XFILLER_136_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6383_ fd._1376_ VGND VGND VPWR VPWR fd._1548_ sky130_fd_sc_hd__clkinvlp_2
XTAP_6180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_261_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_255_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8122_ fd._3428_ fd._3435_ VGND VGND VPWR VPWR fd._3437_ sky130_fd_sc_hd__nor2_1
Xfd._5334_ fd._3580_ fd._0392_ VGND VGND VPWR VPWR fd._0394_ sky130_fd_sc_hd__nand2_1
XFILLER_83_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8053_ fd._3383_ VGND VGND VPWR VPWR fd._3385_ sky130_fd_sc_hd__inv_2
Xfd._5265_ fd._0126_ fd._0130_ VGND VGND VPWR VPWR fd._0319_ sky130_fd_sc_hd__nand2_1
XFILLER_224_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7004_ fd._2025_ VGND VGND VPWR VPWR fd._2231_ sky130_fd_sc_hd__clkinv_2
XFILLER_58_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4216_ fd._1539_ fd._1550_ fd._1220_ VGND VGND VPWR VPWR fd._1561_ sky130_fd_sc_hd__mux2_1
XFILLER_224_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5196_ fd._0070_ fd._0211_ fd._0226_ VGND VGND VPWR VPWR fd._0243_ sky130_fd_sc_hd__and3_1
XFILLER_23_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4147_ fd.b\[12\] fd._0780_ VGND VGND VPWR VPWR fd._0802_ sky130_fd_sc_hd__nand2_1
XFILLER_264_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_264_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4078_ fd.a\[16\] VGND VGND VPWR VPWR fd._0043_ sky130_fd_sc_hd__inv_2
XFILLER_143_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7906_ fd._3043_ fd._3074_ VGND VGND VPWR VPWR fd._3224_ sky130_fd_sc_hd__nor2_1
XFILLER_104_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7837_ fd._2141_ fd._3146_ VGND VGND VPWR VPWR fd._3148_ sky130_fd_sc_hd__or2_1
XFILLER_129_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7768_ fd._2887_ fd._3071_ VGND VGND VPWR VPWR fd._3072_ sky130_fd_sc_hd__xnor2_1
XFILLER_69_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_258_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6719_ fd._1721_ fd._1801_ fd._1917_ VGND VGND VPWR VPWR fd._1918_ sky130_fd_sc_hd__mux2_1
XFILLER_195_1498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7699_ fd._2993_ fd._2994_ fd._2876_ fd._2995_ VGND VGND VPWR VPWR fd._2996_ sky130_fd_sc_hd__o31a_1
XFILLER_132_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_259_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_227_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_265_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_265_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_214_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_230_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_243_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout75 net76 VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_4
XFILLER_11_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_276_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_1671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_284_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5050_ fd._0081_ fd._3979_ fd._0059_ VGND VGND VPWR VPWR fd._0082_ sky130_fd_sc_hd__mux2_1
XFILLER_206_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_283_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_1629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_1517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5952_ fd._1062_ fd._1069_ fd._1072_ fd._1073_ VGND VGND VPWR VPWR fd._1074_ sky130_fd_sc_hd__o211a_1
XFILLER_158_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4903_ fd._3994_ fd._3996_ VGND VGND VPWR VPWR fd._3997_ sky130_fd_sc_hd__xor2_1
XFILLER_220_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5883_ fd._0995_ fd._0996_ fd._0997_ VGND VGND VPWR VPWR fd._0998_ sky130_fd_sc_hd__or3_4
XFILLER_174_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7622_ fd._2909_ fd._2910_ fd._2874_ VGND VGND VPWR VPWR fd._2911_ sky130_fd_sc_hd__mux2_1
Xfd._4834_ fd._3817_ fd._3926_ fd._3927_ VGND VGND VPWR VPWR fd._3928_ sky130_fd_sc_hd__a21oi_1
XFILLER_173_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_259_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4765_ fd._3682_ fd._3699_ VGND VGND VPWR VPWR fd._3859_ sky130_fd_sc_hd__xnor2_1
Xfd._7553_ fd._2831_ fd._2834_ fd._2813_ VGND VGND VPWR VPWR fd._2835_ sky130_fd_sc_hd__mux2_1
XFILLER_118_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_272_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6504_ fd._1319_ fd._1680_ VGND VGND VPWR VPWR fd._1681_ sky130_fd_sc_hd__nor2_1
XFILLER_9_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4696_ fd._3628_ VGND VGND VPWR VPWR fd._3790_ sky130_fd_sc_hd__inv_2
Xfd._7484_ fd._1764_ fd._2577_ fd._2670_ fd._2675_ VGND VGND VPWR VPWR fd._2759_ sky130_fd_sc_hd__o211a_1
XFILLER_142_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_256_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_269_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6435_ fd._1603_ fd._1604_ VGND VGND VPWR VPWR fd._1606_ sky130_fd_sc_hd__and2b_1
XFILLER_68_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_1368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6366_ fd._1321_ fd._1526_ fd._1529_ VGND VGND VPWR VPWR fd._1530_ sky130_fd_sc_hd__mux2_1
XFILLER_3_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_256_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8105_ fd._3800_ fd._3961_ fd._3411_ VGND VGND VPWR VPWR fd._3423_ sky130_fd_sc_hd__mux2_1
XFILLER_231_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._5317_ fd._0180_ VGND VGND VPWR VPWR fd._0376_ sky130_fd_sc_hd__clkinv_2
XFILLER_209_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6297_ fd._0343_ fd._1453_ VGND VGND VPWR VPWR fd._1454_ sky130_fd_sc_hd__nor2_1
XFILLER_3_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5248_ fd._0139_ fd._0299_ fd._0268_ VGND VGND VPWR VPWR fd._0300_ sky130_fd_sc_hd__mux2_1
XFILLER_149_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8036_ fd._3366_ fd._3120_ VGND VGND VPWR VPWR fd._3367_ sky130_fd_sc_hd__xor2_1
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_266_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_251_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5179_ fd._3773_ fd._0221_ VGND VGND VPWR VPWR fd._0224_ sky130_fd_sc_hd__nor2_1
XFILLER_52_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_275_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_1686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_1539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_233_ fd.c\[25\] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_1
XFILLER_230_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_278_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4550_ fd._3277_ fd._3643_ fd._3625_ VGND VGND VPWR VPWR fd._3644_ sky130_fd_sc_hd__mux2_1
XFILLER_139_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_269_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4481_ fd._3574_ VGND VGND VPWR VPWR fd._3575_ sky130_fd_sc_hd__inv_2
XFILLER_133_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_284_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6220_ fd._1178_ fd._1368_ VGND VGND VPWR VPWR fd._1369_ sky130_fd_sc_hd__and2_1
XFILLER_215_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_280_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6151_ fd._1319_ fd._1288_ VGND VGND VPWR VPWR fd._1293_ sky130_fd_sc_hd__and2_1
XFILLER_24_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5102_ fd._0138_ fd._3987_ fd._0060_ VGND VGND VPWR VPWR fd._0139_ sky130_fd_sc_hd__mux2_1
XFILLER_280_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_283_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6082_ fd._1178_ fd._1183_ VGND VGND VPWR VPWR fd._1217_ sky130_fd_sc_hd__and2_1
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_1442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5033_ fd._0015_ fd._0014_ VGND VGND VPWR VPWR fd._0063_ sky130_fd_sc_hd__or2b_1
XFILLER_206_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_283_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_222_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_267_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6984_ fd._2208_ fd._1993_ VGND VGND VPWR VPWR fd._2209_ sky130_fd_sc_hd__xnor2_1
XFILLER_159_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5935_ fd._1042_ fd._0872_ fd._0856_ VGND VGND VPWR VPWR fd._1056_ sky130_fd_sc_hd__o21a_1
XFILLER_119_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5866_ fd._0768_ fd._0867_ VGND VGND VPWR VPWR fd._0980_ sky130_fd_sc_hd__nand2_1
XFILLER_283_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7605_ fd._1494_ fd._2891_ VGND VGND VPWR VPWR fd._2893_ sky130_fd_sc_hd__and2_1
Xfd._4817_ fd._3910_ VGND VGND VPWR VPWR fd._3911_ sky130_fd_sc_hd__clkinv_2
XFILLER_161_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5797_ fd._0683_ fd._0684_ fd._0685_ fd._0687_ VGND VGND VPWR VPWR fd._0904_ sky130_fd_sc_hd__a31o_1
XFILLER_216_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_251_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7536_ fd._2427_ fd._2814_ VGND VGND VPWR VPWR fd._2817_ sky130_fd_sc_hd__and2_1
XFILLER_255_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4748_ fd._3702_ fd._3705_ fd._3709_ VGND VGND VPWR VPWR fd._3842_ sky130_fd_sc_hd__a21o_1
XFILLER_118_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_272_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_257_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7467_ fd._2543_ fd._2740_ fd._2676_ VGND VGND VPWR VPWR fd._2741_ sky130_fd_sc_hd__mux2_1
XFILLER_116_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4679_ fd.b\[21\] VGND VGND VPWR VPWR fd._3773_ sky130_fd_sc_hd__buf_6
XFILLER_233_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6418_ fd._1577_ fd._1586_ VGND VGND VPWR VPWR fd._1587_ sky130_fd_sc_hd__or2b_1
XFILLER_112_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_284_662 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7398_ fd._2623_ fd._2663_ fd._2664_ VGND VGND VPWR VPWR fd._2665_ sky130_fd_sc_hd__a21oi_2
XFILLER_272_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6349_ fd._1507_ fd._1510_ VGND VGND VPWR VPWR fd._1511_ sky130_fd_sc_hd__nand2_1
XFILLER_99_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8019_ fd._3126_ fd._3347_ fd._3239_ VGND VGND VPWR VPWR fd._3348_ sky130_fd_sc_hd__mux2_1
XFILLER_24_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_273_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_8137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_273_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_275_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_262_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_284_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_216_ fd.c\[8\] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_1
XFILLER_141_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5720_ fd._0817_ fd._0818_ VGND VGND VPWR VPWR fd._0819_ sky130_fd_sc_hd__nor2_1
XFILLER_176_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5651_ fd._0742_ VGND VGND VPWR VPWR fd._0743_ sky130_fd_sc_hd__inv_2
XFILLER_143_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._4602_ fd._3695_ fd._3624_ fd._3537_ VGND VGND VPWR VPWR fd._3696_ sky130_fd_sc_hd__o21ai_2
XTAP_8682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5582_ fd._3980_ fd._0665_ VGND VGND VPWR VPWR fd._0667_ sky130_fd_sc_hd__and2_1
XFILLER_112_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7321_ fd._2578_ fd._2394_ VGND VGND VPWR VPWR fd._2580_ sky130_fd_sc_hd__nor2_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4533_ fd._3233_ fd._3584_ fd._3626_ VGND VGND VPWR VPWR fd._3627_ sky130_fd_sc_hd__mux2_1
XTAP_7992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4464_ fd.b\[11\] fd._3553_ fd._3554_ fd._3557_ VGND VGND VPWR VPWR fd._3558_
+ sky130_fd_sc_hd__a31o_1
XFILLER_239_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7252_ fd._2472_ fd._2478_ fd._2480_ fd._2500_ fd._2503_ VGND VGND VPWR VPWR fd._2504_
+ sky130_fd_sc_hd__o221a_2
XFILLER_113_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_254_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6203_ fd._1171_ fd._1228_ fd._1349_ VGND VGND VPWR VPWR fd._1350_ sky130_fd_sc_hd__mux2_1
Xfd._4395_ fd._2177_ fd._3488_ fd._3200_ VGND VGND VPWR VPWR fd._3489_ sky130_fd_sc_hd__mux2_1
Xfd._7183_ fd._2284_ fd._2288_ VGND VGND VPWR VPWR fd._2428_ sky130_fd_sc_hd__nor2_1
XFILLER_113_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_285_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6134_ fd._0541_ fd._1272_ VGND VGND VPWR VPWR fd._1274_ sky130_fd_sc_hd__nor2_1
XFILLER_93_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_263_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6065_ fd._1197_ VGND VGND VPWR VPWR fd._1199_ sky130_fd_sc_hd__clkinv_2
XFILLER_234_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_280_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_278_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5016_ fd._0044_ fd._3952_ VGND VGND VPWR VPWR fd._0045_ sky130_fd_sc_hd__xnor2_1
XFILLER_61_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6967_ fd._1559_ fd._2157_ VGND VGND VPWR VPWR fd._2191_ sky130_fd_sc_hd__or2_1
XFILLER_120_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_1442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5918_ fd._0526_ fd._0988_ VGND VGND VPWR VPWR fd._1037_ sky130_fd_sc_hd__or2_1
XFILLER_175_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6898_ fd._2114_ VGND VGND VPWR VPWR fd._2115_ sky130_fd_sc_hd__buf_6
XFILLER_162_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5849_ fd._0729_ VGND VGND VPWR VPWR fd._0961_ sky130_fd_sc_hd__clkinv_2
XFILLER_162_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_270_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_249_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7519_ fd._2713_ fd._2794_ fd._2796_ fd._2797_ VGND VGND VPWR VPWR fd._2798_ sky130_fd_sc_hd__o211ai_2
XTAP_5319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_268_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_246_1678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_281_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_268_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_251_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_276_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4180_ fd._1143_ VGND VGND VPWR VPWR fd._1165_ sky130_fd_sc_hd__buf_6
XFILLER_263_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_262_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_245_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7870_ fd._2566_ fd._3183_ VGND VGND VPWR VPWR fd._3184_ sky130_fd_sc_hd__and2_1
XFILLER_19_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6821_ fd._1816_ fd._2019_ VGND VGND VPWR VPWR fd._2030_ sky130_fd_sc_hd__nand2_1
XFILLER_15_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_258_1527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6752_ fd._1951_ fd._1953_ VGND VGND VPWR VPWR fd._1954_ sky130_fd_sc_hd__xor2_1
XFILLER_157_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5703_ fd._0785_ fd._0790_ fd._0799_ VGND VGND VPWR VPWR fd._0800_ sky130_fd_sc_hd__o21ai_1
XFILLER_183_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._6683_ fd._1872_ fd._1877_ VGND VGND VPWR VPWR fd._1878_ sky130_fd_sc_hd__nor2_1
XFILLER_144_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_256_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5634_ fd._0656_ fd._0722_ fd._0723_ VGND VGND VPWR VPWR fd._0724_ sky130_fd_sc_hd__a21o_1
XFILLER_125_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5565_ fd._0583_ VGND VGND VPWR VPWR fd._0649_ sky130_fd_sc_hd__clkinv_2
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7304_ fd._2544_ fd._2552_ fd._2558_ fd._2559_ fd._2560_ VGND VGND VPWR VPWR fd._2561_
+ sky130_fd_sc_hd__a311o_1
XFILLER_112_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4516_ fd._3090_ fd._3609_ fd._3222_ VGND VGND VPWR VPWR fd._3610_ sky130_fd_sc_hd__mux2_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_1612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5496_ fd._0369_ fd._0374_ VGND VGND VPWR VPWR fd._0573_ sky130_fd_sc_hd__nand2_1
XFILLER_22_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7235_ fd._2482_ fd._2484_ fd._2423_ VGND VGND VPWR VPWR fd._2486_ sky130_fd_sc_hd__mux2_1
XFILLER_38_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4447_ fd._3531_ fd._3535_ fd._3539_ fd._3540_ VGND VGND VPWR VPWR fd._3541_ sky130_fd_sc_hd__o31a_1
XFILLER_213_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7166_ fd._1661_ fd._2409_ VGND VGND VPWR VPWR fd._2410_ sky130_fd_sc_hd__nor2_1
XFILLER_54_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4378_ fd._2320_ fd._2331_ fd._2342_ fd._2364_ fd._1627_ VGND VGND VPWR VPWR fd._3343_
+ sky130_fd_sc_hd__o311ai_1
XFILLER_199_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6117_ fd._1102_ fd._1255_ VGND VGND VPWR VPWR fd._1256_ sky130_fd_sc_hd__nand2_1
XFILLER_187_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7097_ fd._2326_ fd._2332_ VGND VGND VPWR VPWR fd._2334_ sky130_fd_sc_hd__nand2_1
XFILLER_263_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6048_ fd._1014_ fd._1179_ fd._1030_ VGND VGND VPWR VPWR fd._1180_ sky130_fd_sc_hd__a21oi_1
XFILLER_39_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7999_ fd._3139_ fd._3325_ fd._3240_ VGND VGND VPWR VPWR fd._3326_ sky130_fd_sc_hd__mux2_1
XFILLER_124_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_274_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_254_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_790 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_253_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_268_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5350_ fd._1352_ fd._0400_ VGND VGND VPWR VPWR fd._0412_ sky130_fd_sc_hd__and2_1
XTAP_6373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4301_ fd._1440_ fd._2408_ fd._2485_ fd._2463_ VGND VGND VPWR VPWR fd._2496_ sky130_fd_sc_hd__o31a_1
XFILLER_208_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5281_ fd._3658_ fd._0335_ VGND VGND VPWR VPWR fd._0336_ sky130_fd_sc_hd__nand2_1
XTAP_5683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7020_ fd._2021_ fd._2247_ fd._2248_ VGND VGND VPWR VPWR fd._2249_ sky130_fd_sc_hd__a21oi_2
XTAP_4971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4232_ fd._1660_ fd._1726_ VGND VGND VPWR VPWR fd._1737_ sky130_fd_sc_hd__nand2_1
XFILLER_224_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4163_ fd._0967_ fd.a\[16\] VGND VGND VPWR VPWR fd._0978_ sky130_fd_sc_hd__nor2_1
XFILLER_224_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4094_ fd.b\[4\] VGND VGND VPWR VPWR fd._0219_ sky130_fd_sc_hd__buf_6
XFILLER_189_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_264_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_259_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7922_ fd._3240_ VGND VGND VPWR VPWR fd._3241_ sky130_fd_sc_hd__buf_6
XFILLER_189_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7853_ fd._2959_ fd._3164_ VGND VGND VPWR VPWR fd._3165_ sky130_fd_sc_hd__or2_1
XFILLER_31_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6804_ fd._1656_ fd._2009_ VGND VGND VPWR VPWR fd._2011_ sky130_fd_sc_hd__nor2_1
XFILLER_117_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7784_ fd._3088_ fd._3015_ VGND VGND VPWR VPWR fd._3089_ sky130_fd_sc_hd__nor2_1
XFILLER_69_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4996_ fd._1352_ fd._0022_ VGND VGND VPWR VPWR fd._0023_ sky130_fd_sc_hd__or2_1
XFILLER_195_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6735_ fd._1762_ fd._1773_ VGND VGND VPWR VPWR fd._1936_ sky130_fd_sc_hd__nor2_1
XFILLER_201_1592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6666_ fd._1659_ fd._1662_ fd._1857_ VGND VGND VPWR VPWR fd._1860_ sky130_fd_sc_hd__and3_1
XFILLER_275_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5617_ fd._3905_ fd._0705_ VGND VGND VPWR VPWR fd._0706_ sky130_fd_sc_hd__nor2_1
XFILLER_113_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6597_ fd._1600_ fd._1782_ VGND VGND VPWR VPWR fd._1784_ sky130_fd_sc_hd__nor2_1
XFILLER_224_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_258_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5548_ fd._0262_ fd._0629_ VGND VGND VPWR VPWR fd._0630_ sky130_fd_sc_hd__nand2_1
XFILLER_224_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_273_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8267_ net66 net20 VGND VGND VPWR VPWR fd.b\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5479_ fd._1451_ fd._0553_ VGND VGND VPWR VPWR fd._0554_ sky130_fd_sc_hd__xnor2_1
XFILLER_85_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7218_ fd._2434_ fd._2464_ fd._2466_ VGND VGND VPWR VPWR fd._2467_ sky130_fd_sc_hd__a21oi_1
XFILLER_2_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._8198_ net76 fd.mc\[22\] VGND VGND VPWR VPWR fd.c\[22\] sky130_fd_sc_hd__dfxtp_4
XFILLER_226_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7149_ fd._2152_ fd._2390_ VGND VGND VPWR VPWR fd._2391_ sky130_fd_sc_hd__xnor2_1
XFILLER_226_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_263_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_1430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._4850_ fd._3778_ fd._3943_ fd._3777_ VGND VGND VPWR VPWR fd._3944_ sky130_fd_sc_hd__a21oi_1
XFILLER_51_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_259_1655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_202 VGND VGND VPWR VPWR user_project_wrapper_202/HI la_data_out[80]
+ sky130_fd_sc_hd__conb_1
XFILLER_86_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_213 VGND VGND VPWR VPWR user_project_wrapper_213/HI la_data_out[91]
+ sky130_fd_sc_hd__conb_1
XFILLER_5_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4781_ fd._3689_ fd._3772_ fd._3783_ fd._3785_ VGND VGND VPWR VPWR fd._3875_ sky130_fd_sc_hd__and4_1
XFILLER_182_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_project_wrapper_224 VGND VGND VPWR VPWR user_project_wrapper_224/HI la_data_out[102]
+ sky130_fd_sc_hd__conb_1
XFILLER_127_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_project_wrapper_235 VGND VGND VPWR VPWR user_project_wrapper_235/HI la_data_out[113]
+ sky130_fd_sc_hd__conb_1
XFILLER_181_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_246 VGND VGND VPWR VPWR user_project_wrapper_246/HI la_data_out[124]
+ sky130_fd_sc_hd__conb_1
Xfd._6520_ fd._1690_ fd._1697_ fd._1698_ VGND VGND VPWR VPWR fd._1699_ sky130_fd_sc_hd__a21oi_2
XFILLER_142_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_project_wrapper_257 VGND VGND VPWR VPWR user_project_wrapper_257/HI wbs_dat_o[3]
+ sky130_fd_sc_hd__conb_1
XFILLER_99_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_268 VGND VGND VPWR VPWR user_project_wrapper_268/HI wbs_dat_o[14]
+ sky130_fd_sc_hd__conb_1
XFILLER_29_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_257_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_279 VGND VGND VPWR VPWR user_project_wrapper_279/HI wbs_dat_o[25]
+ sky130_fd_sc_hd__conb_1
XFILLER_194_1680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6451_ fd._1513_ fd._1524_ fd._1522_ VGND VGND VPWR VPWR fd._1623_ sky130_fd_sc_hd__a21boi_1
XFILLER_214_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5402_ fd._3773_ fd._0468_ VGND VGND VPWR VPWR fd._0469_ sky130_fd_sc_hd__nor2_2
XFILLER_150_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._6382_ fd._0928_ fd._1546_ VGND VGND VPWR VPWR fd._1547_ sky130_fd_sc_hd__or2_1
XFILLER_136_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_268_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._8121_ fd._3428_ fd._3435_ VGND VGND VPWR VPWR fd._3436_ sky130_fd_sc_hd__and2_1
XFILLER_256_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5333_ fd._3580_ fd._0392_ VGND VGND VPWR VPWR fd._0393_ sky130_fd_sc_hd__or2_1
XFILLER_0_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_255_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8052_ fd._3356_ fd._3360_ fd._3382_ fd._3383_ VGND VGND VPWR VPWR fd._3384_ sky130_fd_sc_hd__o211a_1
XFILLER_76_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5264_ fd._0312_ fd._0316_ VGND VGND VPWR VPWR fd._0317_ sky130_fd_sc_hd__nor2_1
XFILLER_208_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7003_ fd._2227_ fd._2229_ VGND VGND VPWR VPWR fd._2230_ sky130_fd_sc_hd__nand2_1
Xfd._4215_ fd._0593_ fd._1484_ VGND VGND VPWR VPWR fd._1550_ sky130_fd_sc_hd__xnor2_1
XFILLER_263_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5195_ fd._0062_ fd._0233_ fd._0239_ VGND VGND VPWR VPWR fd._0242_ sky130_fd_sc_hd__a21oi_4
XFILLER_224_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._4146_ fd.b\[12\] fd._0780_ VGND VGND VPWR VPWR fd._0791_ sky130_fd_sc_hd__nor2_1
XFILLER_223_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_260_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4077_ fd.b\[17\] fd._0021_ VGND VGND VPWR VPWR fd._0032_ sky130_fd_sc_hd__nor2_1
XFILLER_225_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7905_ fd._3067_ fd._3080_ fd._3213_ fd._3066_ VGND VGND VPWR VPWR fd._3223_ sky130_fd_sc_hd__a31o_1
XFILLER_137_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_277_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7836_ fd._2141_ fd._3146_ VGND VGND VPWR VPWR fd._3147_ sky130_fd_sc_hd__nand2_1
XFILLER_191_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7767_ fd._2893_ fd._3018_ VGND VGND VPWR VPWR fd._3071_ sky130_fd_sc_hd__nor2_1
Xfd._4979_ fd._0000_ fd._0003_ VGND VGND VPWR VPWR fd._0004_ sky130_fd_sc_hd__nor2_1
XFILLER_144_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6718_ fd._1916_ VGND VGND VPWR VPWR fd._1917_ sky130_fd_sc_hd__buf_6
XFILLER_145_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_254_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7698_ fd._2702_ fd._2876_ VGND VGND VPWR VPWR fd._2995_ sky130_fd_sc_hd__nand2_1
XFILLER_271_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6649_ fd._1837_ fd._1813_ fd._1839_ fd._1840_ VGND VGND VPWR VPWR fd._1841_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_134_1704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_271_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_247_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_274_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_230_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_243_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_265_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout76 net77 VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_6
XFILLER_161_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_254_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_283_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_261_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5951_ fd._0479_ fd._1061_ VGND VGND VPWR VPWR fd._1073_ sky130_fd_sc_hd__nand2_1
XFILLER_119_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4902_ fd._3874_ fd._3995_ VGND VGND VPWR VPWR fd._3996_ sky130_fd_sc_hd__nand2_1
XFILLER_174_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5882_ fd._0886_ fd._0979_ fd._0983_ fd._0873_ VGND VGND VPWR VPWR fd._0997_ sky130_fd_sc_hd__o211a_1
XFILLER_173_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7621_ fd._2785_ fd._2901_ VGND VGND VPWR VPWR fd._2910_ sky130_fd_sc_hd__xnor2_1
Xfd._4833_ fd._1253_ fd._3812_ VGND VGND VPWR VPWR fd._3927_ sky130_fd_sc_hd__nor2_1
XFILLER_127_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7552_ fd._2832_ fd._2833_ VGND VGND VPWR VPWR fd._2834_ sky130_fd_sc_hd__xnor2_1
Xfd._4764_ fd._3669_ fd._3857_ VGND VGND VPWR VPWR fd._3858_ sky130_fd_sc_hd__nand2_1
XFILLER_141_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6503_ fd._1676_ fd._1615_ fd._1678_ fd._1679_ VGND VGND VPWR VPWR fd._1680_ sky130_fd_sc_hd__a22oi_2
XFILLER_272_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_269_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7483_ fd._2751_ fd._2752_ fd._2757_ VGND VGND VPWR VPWR fd._2758_ sky130_fd_sc_hd__and3_1
Xfd._4695_ fd._3759_ fd._3755_ fd._3788_ VGND VGND VPWR VPWR fd._3789_ sky130_fd_sc_hd__mux2_1
XFILLER_233_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6434_ fd._0916_ fd._1602_ VGND VGND VPWR VPWR fd._1604_ sky130_fd_sc_hd__or2_1
XFILLER_151_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_284_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_256_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6365_ fd._1316_ fd._1527_ fd._1314_ VGND VGND VPWR VPWR fd._1529_ sky130_fd_sc_hd__o21ai_1
XFILLER_28_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8104_ fd._3421_ VGND VGND VPWR VPWR fd.mc\[19\] sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5316_ fd._3646_ fd._0369_ fd._0374_ VGND VGND VPWR VPWR fd._0375_ sky130_fd_sc_hd__mux2_1
XFILLER_23_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6296_ fd._1449_ fd._1452_ fd._1422_ VGND VGND VPWR VPWR fd._1453_ sky130_fd_sc_hd__mux2_1
XFILLER_77_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8035_ fd._3119_ fd._3338_ fd._3103_ VGND VGND VPWR VPWR fd._3366_ sky130_fd_sc_hd__a21boi_1
Xfd._5247_ fd._0136_ fd._0298_ VGND VGND VPWR VPWR fd._0299_ sky130_fd_sc_hd__xnor2_1
XFILLER_52_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_266_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5178_ fd._1165_ fd._0222_ VGND VGND VPWR VPWR fd._0223_ sky130_fd_sc_hd__nor2_1
XFILLER_149_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_251_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4129_ fd.b\[8\] fd.a\[8\] VGND VGND VPWR VPWR fd._0604_ sky130_fd_sc_hd__nor2b_1
XFILLER_211_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7819_ fd._3126_ VGND VGND VPWR VPWR fd._3128_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_192_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_259_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_227_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_280_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_232_ fd.c\[24\] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_1
XFILLER_211_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_266_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4480_ fd._3569_ fd._3573_ VGND VGND VPWR VPWR fd._3574_ sky130_fd_sc_hd__nand2_1
XFILLER_6_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_1667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6150_ fd._1291_ VGND VGND VPWR VPWR fd._1292_ sky130_fd_sc_hd__clkinv_4
XFILLER_20_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5101_ fd._3990_ fd._0137_ VGND VGND VPWR VPWR fd._0138_ sky130_fd_sc_hd__xnor2_1
XFILLER_19_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6081_ fd._1196_ fd._1205_ fd._1213_ fd._1214_ fd._1215_ VGND VGND VPWR VPWR fd._1216_
+ sky130_fd_sc_hd__a311o_1
XFILLER_34_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_283_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5032_ fd._3963_ fd._0042_ fd._0061_ VGND VGND VPWR VPWR fd._0062_ sky130_fd_sc_hd__mux2_4
XFILLER_185_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6983_ fd._1996_ fd._2207_ fd._1931_ VGND VGND VPWR VPWR fd._2208_ sky130_fd_sc_hd__o21a_1
XFILLER_144_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5934_ fd._0855_ fd._1042_ fd._1047_ VGND VGND VPWR VPWR fd._1054_ sky130_fd_sc_hd__a21oi_1
XFILLER_140_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5865_ fd._0970_ fd._0973_ fd._0975_ fd._0977_ VGND VGND VPWR VPWR fd._0979_ sky130_fd_sc_hd__o211a_1
XFILLER_179_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7604_ fd._2808_ fd._2890_ fd._2875_ VGND VGND VPWR VPWR fd._2891_ sky130_fd_sc_hd__mux2_1
XFILLER_283_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4816_ fd._3909_ fd._3712_ VGND VGND VPWR VPWR fd._3910_ sky130_fd_sc_hd__xnor2_1
XFILLER_196_1583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5796_ fd._0716_ fd._0902_ VGND VGND VPWR VPWR fd._0903_ sky130_fd_sc_hd__or2_1
XFILLER_143_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7535_ fd._2427_ fd._2814_ VGND VGND VPWR VPWR fd._2816_ sky130_fd_sc_hd__nor2_1
Xfd._4747_ fd._3839_ fd._3840_ VGND VGND VPWR VPWR fd._3841_ sky130_fd_sc_hd__nor2_1
XFILLER_142_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_272_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_269_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7466_ fd._2544_ fd._2739_ VGND VGND VPWR VPWR fd._2740_ sky130_fd_sc_hd__xnor2_1
Xfd._4678_ fd._3763_ fd._3767_ fd._3770_ fd._3771_ VGND VGND VPWR VPWR fd._3772_ sky130_fd_sc_hd__a211oi_2
XFILLER_257_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6417_ fd._1585_ fd._1399_ VGND VGND VPWR VPWR fd._1586_ sky130_fd_sc_hd__nand2_1
XFILLER_68_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7397_ fd._2475_ fd._2623_ VGND VGND VPWR VPWR fd._2664_ sky130_fd_sc_hd__nor2_1
XFILLER_9_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_284_674 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6348_ fd._1326_ fd._1509_ fd._1423_ VGND VGND VPWR VPWR fd._1510_ sky130_fd_sc_hd__mux2_1
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6279_ fd._1431_ fd._1433_ VGND VGND VPWR VPWR fd._1434_ sky130_fd_sc_hd__nand2_1
XFILLER_37_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._8018_ fd._3344_ fd._3346_ VGND VGND VPWR VPWR fd._3347_ sky130_fd_sc_hd__xnor2_1
XFILLER_225_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_273_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_275_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_1484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_284_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_1662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_1657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_215_ fd.c\[7\] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_1
XFILLER_50_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_258_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5650_ fd._0576_ fd._0741_ fd._0651_ VGND VGND VPWR VPWR fd._0742_ sky130_fd_sc_hd__mux2_1
XFILLER_256_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4601_ fd._3536_ VGND VGND VPWR VPWR fd._3695_ sky130_fd_sc_hd__buf_6
XTAP_8672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5581_ fd._0662_ fd._0665_ VGND VGND VPWR VPWR fd._0666_ sky130_fd_sc_hd__nor2_1
XTAP_8694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7320_ fd._2578_ fd._2394_ VGND VGND VPWR VPWR fd._2579_ sky130_fd_sc_hd__and2_1
XFILLER_139_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4532_ fd._3625_ VGND VGND VPWR VPWR fd._3626_ sky130_fd_sc_hd__buf_6
XTAP_7971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_1617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7251_ fd._2502_ fd._2501_ fd._2239_ VGND VGND VPWR VPWR fd._2503_ sky130_fd_sc_hd__mux2_1
Xfd._4463_ fd._1594_ fd._3556_ fd._3211_ VGND VGND VPWR VPWR fd._3557_ sky130_fd_sc_hd__mux2_1
XFILLER_6_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6202_ fd._1340_ fd._1348_ VGND VGND VPWR VPWR fd._1349_ sky130_fd_sc_hd__nand2_4
XFILLER_120_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7182_ fd._1431_ VGND VGND VPWR VPWR fd._2427_ sky130_fd_sc_hd__buf_6
XFILLER_66_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._4394_ fd._3387_ fd._3479_ VGND VGND VPWR VPWR fd._3488_ sky130_fd_sc_hd__or2b_1
XFILLER_4_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_280_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6133_ fd._0541_ fd._1272_ VGND VGND VPWR VPWR fd._1273_ sky130_fd_sc_hd__nand2_1
XFILLER_207_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6064_ fd._0985_ fd._1021_ fd._1024_ VGND VGND VPWR VPWR fd._1197_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_267_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_1568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5015_ fd._3937_ fd._3942_ VGND VGND VPWR VPWR fd._0044_ sky130_fd_sc_hd__nand2_1
XFILLER_222_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6966_ fd._2142_ fd._2164_ VGND VGND VPWR VPWR fd._2190_ sky130_fd_sc_hd__nand2_1
XFILLER_119_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5917_ fd._0526_ fd._0988_ VGND VGND VPWR VPWR fd._1036_ sky130_fd_sc_hd__nand2_1
XFILLER_190_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6897_ fd._2033_ fd._2048_ fd._2113_ VGND VGND VPWR VPWR fd._2114_ sky130_fd_sc_hd__or3_1
XFILLER_135_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5848_ fd._0897_ fd._0953_ fd._0959_ fd._0895_ VGND VGND VPWR VPWR fd._0960_ sky130_fd_sc_hd__a31oi_2
XFILLER_66_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_1664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_1498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5779_ fd._0594_ fd._0883_ VGND VGND VPWR VPWR fd._0884_ sky130_fd_sc_hd__nor2_1
XFILLER_130_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7518_ fd._2710_ VGND VGND VPWR VPWR fd._2797_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_115_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_257_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7449_ fd._1219_ fd._2522_ VGND VGND VPWR VPWR fd._2721_ sky130_fd_sc_hd__or2_1
XFILLER_131_1504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_257_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_272_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_281_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_273_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_283_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_262_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_251_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_284_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1590 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6820_ fd._1815_ fd._2028_ VGND VGND VPWR VPWR fd._2029_ sky130_fd_sc_hd__xnor2_1
XFILLER_141_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6751_ fd._1762_ fd._1952_ VGND VGND VPWR VPWR fd._1953_ sky130_fd_sc_hd__nor2_1
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5702_ fd._0797_ fd._0798_ fd._0455_ VGND VGND VPWR VPWR fd._0799_ sky130_fd_sc_hd__mux2_1
XFILLER_176_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6682_ fd._1874_ fd._1875_ fd._1720_ fd._1876_ VGND VGND VPWR VPWR fd._1877_ sky130_fd_sc_hd__a31o_1
XTAP_9170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_1640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_9181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5633_ fd._3917_ fd._0661_ fd._0721_ VGND VGND VPWR VPWR fd._0723_ sky130_fd_sc_hd__and3_1
XFILLER_252_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_252_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5564_ fd._0643_ fd._0646_ VGND VGND VPWR VPWR fd._0647_ sky130_fd_sc_hd__xnor2_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_1559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7303_ fd._1559_ fd._2537_ VGND VGND VPWR VPWR fd._2560_ sky130_fd_sc_hd__nor2_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4515_ fd._3607_ fd._3608_ VGND VGND VPWR VPWR fd._3609_ sky130_fd_sc_hd__xnor2_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5495_ fd._3646_ fd._0569_ fd._0570_ VGND VGND VPWR VPWR fd._0572_ sky130_fd_sc_hd__a21o_1
XFILLER_112_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7234_ fd._2291_ fd._2483_ VGND VGND VPWR VPWR fd._2484_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4446_ fd.b\[3\] fd._3530_ VGND VGND VPWR VPWR fd._3540_ sky130_fd_sc_hd__or2_1
XFILLER_113_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_281_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_269_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7165_ fd._2218_ fd._2407_ fd._2323_ VGND VGND VPWR VPWR fd._2409_ sky130_fd_sc_hd__mux2_1
XFILLER_113_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4377_ fd._1297_ fd._3277_ fd._3321_ VGND VGND VPWR VPWR fd._3332_ sky130_fd_sc_hd__a21oi_1
XFILLER_226_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6116_ fd._1082_ fd._1254_ fd._1223_ VGND VGND VPWR VPWR fd._1255_ sky130_fd_sc_hd__mux2_1
XFILLER_187_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._7096_ fd._2326_ fd._2332_ VGND VGND VPWR VPWR fd._2333_ sky130_fd_sc_hd__or2_1
XFILLER_39_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_263_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6047_ fd._1020_ fd._1029_ VGND VGND VPWR VPWR fd._1179_ sky130_fd_sc_hd__and2_1
XFILLER_250_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._7998_ fd._3323_ fd._3324_ VGND VGND VPWR VPWR fd._3325_ sky130_fd_sc_hd__xnor2_1
XFILLER_120_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6949_ fd._1975_ fd._2168_ fd._2169_ VGND VGND VPWR VPWR fd._2171_ sky130_fd_sc_hd__a21oi_1
XFILLER_162_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_252_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_249_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_264_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_270_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_281_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_257_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4300_ fd._2463_ fd._2474_ VGND VGND VPWR VPWR fd._2485_ sky130_fd_sc_hd__nand2_1
XFILLER_267_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5280_ fd._0332_ fd._0269_ fd._0333_ fd._0334_ VGND VGND VPWR VPWR fd._0335_ sky130_fd_sc_hd__a31o_1
XTAP_5673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._4231_ fd._0230_ fd._1649_ VGND VGND VPWR VPWR fd._1726_ sky130_fd_sc_hd__or2_1
XFILLER_169_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4162_ fd.b\[16\] VGND VGND VPWR VPWR fd._0967_ sky130_fd_sc_hd__clkinv_4
XFILLER_263_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4093_ fd._0186_ fd._0197_ VGND VGND VPWR VPWR fd._0208_ sky130_fd_sc_hd__or2_1
XFILLER_232_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_1685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_225_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7921_ fd._3239_ VGND VGND VPWR VPWR fd._3240_ sky130_fd_sc_hd__buf_6
XFILLER_149_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._7852_ fd._2377_ fd._1970_ fd._2876_ VGND VGND VPWR VPWR fd._3164_ sky130_fd_sc_hd__and3_1
XFILLER_121_1503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6803_ fd._1656_ fd._2009_ VGND VGND VPWR VPWR fd._2010_ sky130_fd_sc_hd__nand2_1
XFILLER_157_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7783_ fd._1685_ fd._3012_ VGND VGND VPWR VPWR fd._3088_ sky130_fd_sc_hd__nor2_1
XFILLER_89_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4995_ fd._3807_ fd._0020_ fd._3961_ VGND VGND VPWR VPWR fd._0022_ sky130_fd_sc_hd__mux2_1
XFILLER_144_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_258_1336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6734_ fd._1751_ fd._1755_ VGND VGND VPWR VPWR fd._1934_ sky130_fd_sc_hd__nand2_1
XFILLER_258_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_275_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6665_ fd._1659_ fd._1662_ fd._1857_ VGND VGND VPWR VPWR fd._1859_ sky130_fd_sc_hd__a21oi_1
XFILLER_208_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5616_ fd._0495_ fd._0704_ fd._0614_ VGND VGND VPWR VPWR fd._0705_ sky130_fd_sc_hd__mux2_1
XFILLER_158_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_256_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6596_ fd._1600_ fd._1782_ VGND VGND VPWR VPWR fd._1783_ sky130_fd_sc_hd__and2_1
XFILLER_99_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5547_ fd._0442_ fd._0628_ fd._0613_ VGND VGND VPWR VPWR fd._0629_ sky130_fd_sc_hd__mux2_1
XFILLER_119_1498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8266_ net66 net19 VGND VGND VPWR VPWR fd.b\[26\] sky130_fd_sc_hd__dfxtp_1
Xfd._5478_ fd._0359_ fd._0552_ fd._0452_ VGND VGND VPWR VPWR fd._0553_ sky130_fd_sc_hd__mux2_1
XFILLER_41_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7217_ fd._2465_ fd._2424_ VGND VGND VPWR VPWR fd._2466_ sky130_fd_sc_hd__nor2_1
XFILLER_82_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4429_ fd._1946_ fd._1957_ VGND VGND VPWR VPWR fd._3523_ sky130_fd_sc_hd__or2_1
XFILLER_187_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8197_ net69 fd.mc\[21\] VGND VGND VPWR VPWR fd.c\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_269_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_270_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7148_ fd._2158_ fd._2192_ VGND VGND VPWR VPWR fd._2390_ sky130_fd_sc_hd__nor2_1
XFILLER_54_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7079_ fd._2304_ fd._2313_ VGND VGND VPWR VPWR fd._2314_ sky130_fd_sc_hd__nand2_1
XFILLER_228_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_276_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_250_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_project_wrapper_203 VGND VGND VPWR VPWR user_project_wrapper_203/HI la_data_out[81]
+ sky130_fd_sc_hd__conb_1
Xfd._4780_ fd._3869_ fd._3873_ VGND VGND VPWR VPWR fd._3874_ sky130_fd_sc_hd__nand2_1
XFILLER_126_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_214 VGND VGND VPWR VPWR user_project_wrapper_214/HI la_data_out[92]
+ sky130_fd_sc_hd__conb_1
XFILLER_86_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_project_wrapper_225 VGND VGND VPWR VPWR user_project_wrapper_225/HI la_data_out[103]
+ sky130_fd_sc_hd__conb_1
XFILLER_5_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_236 VGND VGND VPWR VPWR user_project_wrapper_236/HI la_data_out[114]
+ sky130_fd_sc_hd__conb_1
XFILLER_181_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_247 VGND VGND VPWR VPWR user_project_wrapper_247/HI la_data_out[125]
+ sky130_fd_sc_hd__conb_1
XFILLER_4_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_258 VGND VGND VPWR VPWR user_project_wrapper_258/HI wbs_dat_o[4]
+ sky130_fd_sc_hd__conb_1
XFILLER_68_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_269 VGND VGND VPWR VPWR user_project_wrapper_269/HI wbs_dat_o[15]
+ sky130_fd_sc_hd__conb_1
XFILLER_5_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6450_ fd._0786_ fd._1621_ VGND VGND VPWR VPWR fd._1622_ sky130_fd_sc_hd__nor2_1
XFILLER_194_1692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5401_ fd._0408_ fd._0467_ fd._0453_ VGND VGND VPWR VPWR fd._0468_ sky130_fd_sc_hd__mux2_1
XFILLER_214_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._6381_ fd._1368_ fd._1545_ fd._1533_ VGND VGND VPWR VPWR fd._1546_ sky130_fd_sc_hd__mux2_1
XTAP_6160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._8120_ fd._3425_ fd._3434_ VGND VGND VPWR VPWR fd._3435_ sky130_fd_sc_hd__xnor2_1
XFILLER_255_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5332_ fd._0073_ fd._0391_ fd._0270_ VGND VGND VPWR VPWR fd._0392_ sky130_fd_sc_hd__mux2_1
XTAP_6193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._8051_ fd._1286_ fd._3380_ fd._3368_ fd._2055_ VGND VGND VPWR VPWR fd._3383_ sky130_fd_sc_hd__o22a_1
XFILLER_114_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5263_ fd._0313_ fd._0315_ fd._0268_ VGND VGND VPWR VPWR fd._0316_ sky130_fd_sc_hd__mux2_1
XFILLER_36_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7002_ fd._2124_ fd._2228_ fd._2226_ VGND VGND VPWR VPWR fd._2229_ sky130_fd_sc_hd__o21ai_1
XFILLER_75_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4214_ fd.a\[10\] VGND VGND VPWR VPWR fd._1539_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_224_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5194_ fd._0062_ fd._0235_ fd._0236_ fd._0239_ VGND VGND VPWR VPWR fd._0240_ sky130_fd_sc_hd__a211o_1
XFILLER_223_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4145_ fd.a\[12\] VGND VGND VPWR VPWR fd._0780_ sky130_fd_sc_hd__inv_2
XFILLER_127_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4076_ fd.a\[17\] VGND VGND VPWR VPWR fd._0021_ sky130_fd_sc_hd__inv_2
XFILLER_182_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7904_ fd._2863_ fd._3220_ VGND VGND VPWR VPWR fd._3221_ sky130_fd_sc_hd__nand2_1
XFILLER_143_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7835_ fd._2935_ fd._3144_ fd._3075_ VGND VGND VPWR VPWR fd._3146_ sky130_fd_sc_hd__mux2_1
XFILLER_125_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_1412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4978_ fd._3820_ fd._0002_ fd._3960_ VGND VGND VPWR VPWR fd._0003_ sky130_fd_sc_hd__mux2_1
Xfd._7766_ fd._2884_ VGND VGND VPWR VPWR fd._3070_ sky130_fd_sc_hd__clkinv_2
XFILLER_69_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._6717_ fd._1821_ fd._1835_ fd._1915_ VGND VGND VPWR VPWR fd._1916_ sky130_fd_sc_hd__nand3_2
XFILLER_105_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._7697_ fd._2800_ fd._2707_ fd._2798_ VGND VGND VPWR VPWR fd._2994_ sky130_fd_sc_hd__and3_1
XFILLER_144_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6648_ fd._1699_ fd._1838_ VGND VGND VPWR VPWR fd._1840_ sky130_fd_sc_hd__nor2_1
XFILLER_232_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._6579_ fd._3695_ VGND VGND VPWR VPWR fd._1764_ sky130_fd_sc_hd__buf_6
XFILLER_150_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8249_ net73 net32 VGND VGND VPWR VPWR fd.b\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_100_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout66 net67 VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_4
XFILLER_168_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout77 net33 VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__buf_8
XFILLER_278_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_250_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_265_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_261_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_265_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5950_ fd._1048_ fd._1071_ VGND VGND VPWR VPWR fd._1072_ sky130_fd_sc_hd__nor2_1
XFILLER_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4901_ fd._3869_ fd._3873_ VGND VGND VPWR VPWR fd._3995_ sky130_fd_sc_hd__or2_1
XFILLER_224_1390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5881_ fd._0874_ VGND VGND VPWR VPWR fd._0996_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_158_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4832_ fd._3821_ fd._3923_ fd._3925_ VGND VGND VPWR VPWR fd._3926_ sky130_fd_sc_hd__a21o_1
Xfd._7620_ fd._2724_ VGND VGND VPWR VPWR fd._2909_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_31_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4763_ fd._3856_ fd._3673_ fd._3787_ VGND VGND VPWR VPWR fd._3857_ sky130_fd_sc_hd__mux2_1
Xfd._7551_ fd._2641_ fd._2655_ VGND VGND VPWR VPWR fd._2833_ sky130_fd_sc_hd__nand2_1
XFILLER_5_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6502_ fd._1675_ fd._1677_ VGND VGND VPWR VPWR fd._1679_ sky130_fd_sc_hd__nand2_1
XFILLER_142_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7482_ fd._2670_ fd._2675_ fd._2755_ fd._2756_ VGND VGND VPWR VPWR fd._2757_ sky130_fd_sc_hd__a211o_1
XFILLER_272_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4694_ fd._3787_ VGND VGND VPWR VPWR fd._3788_ sky130_fd_sc_hd__buf_6
XFILLER_272_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_253_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6433_ fd._1600_ fd._1602_ VGND VGND VPWR VPWR fd._1603_ sky130_fd_sc_hd__and2_1
XFILLER_9_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_268_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_269_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_256_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6364_ fd._1516_ VGND VGND VPWR VPWR fd._1527_ sky130_fd_sc_hd__inv_2
XFILLER_68_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8103_ fd._3961_ fd._0061_ fd._3411_ VGND VGND VPWR VPWR fd._3421_ sky130_fd_sc_hd__mux2_1
Xfd._5315_ fd._3646_ fd._0372_ VGND VGND VPWR VPWR fd._0374_ sky130_fd_sc_hd__xnor2_1
XFILLER_42_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6295_ fd._1450_ fd._1265_ VGND VGND VPWR VPWR fd._1452_ sky130_fd_sc_hd__xnor2_1
XFILLER_37_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8034_ fd._2465_ fd._3363_ VGND VGND VPWR VPWR fd._3364_ sky130_fd_sc_hd__nand2_1
Xfd._5246_ fd._0297_ fd._0140_ VGND VGND VPWR VPWR fd._0298_ sky130_fd_sc_hd__nor2_1
XFILLER_225_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5177_ fd._0221_ VGND VGND VPWR VPWR fd._0222_ sky130_fd_sc_hd__inv_2
XFILLER_224_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4128_ fd._0571_ fd._0582_ VGND VGND VPWR VPWR fd._0593_ sky130_fd_sc_hd__nor2_1
XFILLER_225_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7818_ fd._1656_ fd._3126_ VGND VGND VPWR VPWR fd._3127_ sky130_fd_sc_hd__nand2_1
XTAP_8309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_273_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_246_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7749_ fd._3050_ VGND VGND VPWR VPWR fd._3051_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_106_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_259_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_231_ fd.c\[23\] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_1
XFILLER_230_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_276_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_285_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_277_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_253_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5100_ fd._3993_ fd._4018_ VGND VGND VPWR VPWR fd._0137_ sky130_fd_sc_hd__or2_1
XFILLER_219_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_283_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6080_ fd._0807_ fd._1188_ VGND VGND VPWR VPWR fd._1215_ sky130_fd_sc_hd__nor2_1
XFILLER_74_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5031_ fd._0060_ VGND VGND VPWR VPWR fd._0061_ sky130_fd_sc_hd__inv_2
XFILLER_65_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6982_ fd._2197_ VGND VGND VPWR VPWR fd._2207_ sky130_fd_sc_hd__inv_2
XFILLER_261_1387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5933_ fd._0786_ fd._1043_ VGND VGND VPWR VPWR fd._1053_ sky130_fd_sc_hd__nand2_1
XFILLER_119_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5864_ fd._0976_ fd._0878_ VGND VGND VPWR VPWR fd._0977_ sky130_fd_sc_hd__nor2_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._7603_ fd._2888_ fd._2889_ VGND VGND VPWR VPWR fd._2890_ sky130_fd_sc_hd__xnor2_1
XFILLER_127_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4815_ fd._3654_ fd._3900_ fd._3713_ VGND VGND VPWR VPWR fd._3909_ sky130_fd_sc_hd__o21a_1
XFILLER_143_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5795_ fd._0711_ fd._0900_ fd._0848_ VGND VGND VPWR VPWR fd._0902_ sky130_fd_sc_hd__mux2_1
XFILLER_6_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4746_ fd._3833_ fd._3838_ VGND VGND VPWR VPWR fd._3840_ sky130_fd_sc_hd__nor2_1
XFILLER_143_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7534_ fd._2651_ fd._2812_ fd._2813_ VGND VGND VPWR VPWR fd._2814_ sky130_fd_sc_hd__mux2_1
XFILLER_255_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4677_ fd._3617_ fd._3626_ fd._3769_ VGND VGND VPWR VPWR fd._3771_ sky130_fd_sc_hd__and3_1
XFILLER_216_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7465_ fd._2552_ fd._2558_ VGND VGND VPWR VPWR fd._2739_ sky130_fd_sc_hd__and2_1
XFILLER_229_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6416_ fd._0632_ VGND VGND VPWR VPWR fd._1585_ sky130_fd_sc_hd__buf_6
XFILLER_151_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7396_ fd._2662_ fd._2479_ VGND VGND VPWR VPWR fd._2663_ sky130_fd_sc_hd__xor2_1
XFILLER_64_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_256_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6347_ fd._1508_ fd._1329_ VGND VGND VPWR VPWR fd._1509_ sky130_fd_sc_hd__xnor2_1
XFILLER_151_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput1 io_in[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_4
XFILLER_284_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6278_ fd._1233_ fd._1432_ VGND VGND VPWR VPWR fd._1433_ sky130_fd_sc_hd__xnor2_1
XFILLER_209_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5229_ fd._0277_ fd._0278_ VGND VGND VPWR VPWR fd._0279_ sky130_fd_sc_hd__nand2_1
Xfd._8017_ fd._3127_ fd._3345_ VGND VGND VPWR VPWR fd._3346_ sky130_fd_sc_hd__and2_1
XFILLER_240_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_262_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_273_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_273_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_251_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_267_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_255_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_251_1534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_259_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_262_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_214_ fd.c\[6\] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_1
XFILLER_223_1669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4600_ fd._3688_ fd._3693_ VGND VGND VPWR VPWR fd._3694_ sky130_fd_sc_hd__nand2_1
XFILLER_87_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5580_ fd._0530_ fd._0664_ fd._0614_ VGND VGND VPWR VPWR fd._0665_ sky130_fd_sc_hd__mux2_1
XFILLER_125_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4531_ fd._3624_ VGND VGND VPWR VPWR fd._3625_ sky130_fd_sc_hd__buf_6
XTAP_7961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7250_ fd._2249_ fd._2501_ VGND VGND VPWR VPWR fd._2502_ sky130_fd_sc_hd__nand2_1
Xfd._4462_ fd._2320_ fd._2342_ VGND VGND VPWR VPWR fd._3556_ sky130_fd_sc_hd__xnor2_1
XFILLER_61_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._6201_ fd._1343_ fd._1344_ fd._1345_ fd._1347_ VGND VGND VPWR VPWR fd._1348_ sky130_fd_sc_hd__o211a_2
XFILLER_117_1596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7181_ fd._0131_ fd._2425_ VGND VGND VPWR VPWR fd._2426_ sky130_fd_sc_hd__nor2_1
XFILLER_120_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4393_ fd._2144_ fd._2221_ VGND VGND VPWR VPWR fd._3479_ sky130_fd_sc_hd__nand2_1
XFILLER_238_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6132_ fd._1100_ fd._1271_ fd._1223_ VGND VGND VPWR VPWR fd._1272_ sky130_fd_sc_hd__mux2_2
XFILLER_187_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_280_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6063_ fd._0427_ fd._1195_ VGND VGND VPWR VPWR fd._1196_ sky130_fd_sc_hd__xnor2_1
XFILLER_146_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_280_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5014_ fd._0038_ fd._0041_ VGND VGND VPWR VPWR fd._0042_ sky130_fd_sc_hd__xor2_1
XFILLER_61_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_261_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6965_ fd._1958_ fd._2173_ fd._2184_ fd._2187_ VGND VGND VPWR VPWR fd._2189_ sky130_fd_sc_hd__o211a_1
XFILLER_124_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5916_ fd._1001_ fd._1034_ VGND VGND VPWR VPWR fd._1035_ sky130_fd_sc_hd__nand2_1
XFILLER_175_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6896_ fd._2063_ fd._2108_ fd._2109_ fd._2110_ fd._2112_ VGND VGND VPWR VPWR fd._2113_
+ sky130_fd_sc_hd__o2111a_1
XFILLER_190_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5847_ fd._3917_ fd._0903_ fd._0952_ fd._0958_ VGND VGND VPWR VPWR fd._0959_ sky130_fd_sc_hd__a31o_1
XFILLER_179_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5778_ fd._0652_ fd._0882_ fd._0849_ VGND VGND VPWR VPWR fd._0883_ sky130_fd_sc_hd__mux2_1
XFILLER_157_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_274_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7517_ fd._2707_ fd._2795_ VGND VGND VPWR VPWR fd._2796_ sky130_fd_sc_hd__and2_1
Xfd._4729_ fd._3821_ fd._3822_ VGND VGND VPWR VPWR fd._3823_ sky130_fd_sc_hd__nand2_1
XFILLER_170_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_233_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7448_ fd._2532_ fd._2538_ fd._2561_ fd._2564_ VGND VGND VPWR VPWR fd._2720_ sky130_fd_sc_hd__a31o_1
XTAP_4609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7379_ fd._2458_ fd._2643_ VGND VGND VPWR VPWR fd._2644_ sky130_fd_sc_hd__xnor2_1
XFILLER_29_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_272_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_281_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_279_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_268_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_1388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_257_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_1629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_284_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_280_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_262_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6750_ fd._1015_ fd._1761_ VGND VGND VPWR VPWR fd._1952_ sky130_fd_sc_hd__nor2_1
XFILLER_157_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5701_ fd._0464_ fd._0797_ VGND VGND VPWR VPWR fd._0798_ sky130_fd_sc_hd__or2b_1
XFILLER_32_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._6681_ fd._1654_ fd._1720_ VGND VGND VPWR VPWR fd._1876_ sky130_fd_sc_hd__nor2_1
XFILLER_171_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5632_ fd._0661_ fd._0721_ fd._3917_ VGND VGND VPWR VPWR fd._0722_ sky130_fd_sc_hd__a21o_1
XTAP_8470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_8481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5563_ fd._0644_ fd._0645_ VGND VGND VPWR VPWR fd._0646_ sky130_fd_sc_hd__nor2_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7302_ fd._1751_ fd._2543_ VGND VGND VPWR VPWR fd._2559_ sky130_fd_sc_hd__nor2_1
XFILLER_112_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4514_ fd._3123_ fd._3112_ VGND VGND VPWR VPWR fd._3608_ sky130_fd_sc_hd__and2b_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_267_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5494_ fd._0564_ fd._0568_ VGND VGND VPWR VPWR fd._0570_ sky130_fd_sc_hd__and2_1
XFILLER_6_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4445_ fd.b\[2\] fd._3534_ fd._3538_ VGND VGND VPWR VPWR fd._3539_ sky130_fd_sc_hd__o21ba_1
Xfd._7233_ fd._2296_ fd._2295_ VGND VGND VPWR VPWR fd._2483_ sky130_fd_sc_hd__or2b_1
XFILLER_269_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_254_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4376_ fd.b\[15\] fd._3277_ fd._3310_ fd.b\[14\] VGND VGND VPWR VPWR fd._3321_
+ sky130_fd_sc_hd__o22a_1
Xfd._7164_ fd._2405_ fd._2406_ VGND VGND VPWR VPWR fd._2407_ sky130_fd_sc_hd__xnor2_1
XFILLER_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6115_ fd._1252_ fd._1094_ VGND VGND VPWR VPWR fd._1254_ sky130_fd_sc_hd__xnor2_1
XFILLER_241_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7095_ fd._2327_ fd._2330_ fd._2323_ VGND VGND VPWR VPWR fd._2332_ sky130_fd_sc_hd__mux2_1
XFILLER_78_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_263_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6046_ fd._1341_ VGND VGND VPWR VPWR fd._1178_ sky130_fd_sc_hd__buf_6
XFILLER_165_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_263_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7997_ fd._3140_ fd._3179_ VGND VGND VPWR VPWR fd._3324_ sky130_fd_sc_hd__or2b_1
XFILLER_175_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6948_ fd._1975_ fd._2168_ fd._2169_ VGND VGND VPWR VPWR fd._2170_ sky130_fd_sc_hd__and3_1
XFILLER_135_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6879_ fd._2093_ fd._2087_ VGND VGND VPWR VPWR fd._2094_ sky130_fd_sc_hd__nand2_1
XFILLER_11_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_249_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_252_1695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_273_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_272_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_1499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_268_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_267_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4230_ fd.a\[4\] VGND VGND VPWR VPWR fd._1715_ sky130_fd_sc_hd__clkinv_2
XFILLER_235_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4161_ fd._0824_ fd._0912_ fd._0934_ fd._0945_ VGND VGND VPWR VPWR fd._0956_ sky130_fd_sc_hd__o211a_1
XFILLER_251_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_1620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_223_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4092_ fd.b\[7\] fd.a\[7\] VGND VGND VPWR VPWR fd._0197_ sky130_fd_sc_hd__xor2_1
XFILLER_1_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7920_ fd._3221_ fd._3230_ fd._3235_ fd._3238_ VGND VGND VPWR VPWR fd._3239_ sky130_fd_sc_hd__a31o_4
XFILLER_147_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._7851_ fd._2751_ fd._3162_ VGND VGND VPWR VPWR fd._3163_ sky130_fd_sc_hd__or2_1
XPHY_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6802_ fd._2007_ fd._1969_ fd._2008_ VGND VGND VPWR VPWR fd._2009_ sky130_fd_sc_hd__o21ai_1
XFILLER_30_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7782_ fd._2427_ fd._3086_ VGND VGND VPWR VPWR fd._3087_ sky130_fd_sc_hd__nor2_1
XFILLER_117_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4994_ fd._0019_ VGND VGND VPWR VPWR fd._0020_ sky130_fd_sc_hd__clkinv_2
XFILLER_160_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6733_ fd._1925_ fd._1931_ fd._1932_ VGND VGND VPWR VPWR fd._1933_ sky130_fd_sc_hd__a21o_1
XFILLER_258_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_275_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_1624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6664_ fd._1667_ fd._1665_ VGND VGND VPWR VPWR fd._1857_ sky130_fd_sc_hd__or2b_1
XFILLER_172_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_256_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5615_ fd._0701_ fd._0702_ VGND VGND VPWR VPWR fd._0704_ sky130_fd_sc_hd__or2_1
XFILLER_154_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_271_1548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_217_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6595_ fd._1540_ fd._1780_ fd._1719_ VGND VGND VPWR VPWR fd._1782_ sky130_fd_sc_hd__mux2_1
XFILLER_112_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5546_ fd._0624_ fd._0627_ VGND VGND VPWR VPWR fd._0628_ sky130_fd_sc_hd__xnor2_1
XFILLER_112_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_255_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8265_ net67 net18 VGND VGND VPWR VPWR fd.b\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_224_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5477_ fd._0350_ fd._0551_ VGND VGND VPWR VPWR fd._0552_ sky130_fd_sc_hd__xnor2_1
XFILLER_67_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7216_ fd._1304_ VGND VGND VPWR VPWR fd._2465_ sky130_fd_sc_hd__buf_6
XFILLER_269_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_255_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4428_ fd._3520_ fd._3521_ VGND VGND VPWR VPWR fd._3522_ sky130_fd_sc_hd__nand2_1
XFILLER_113_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._8196_ net69 fd.mc\[20\] VGND VGND VPWR VPWR fd.c\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_226_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1690 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_281_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4359_ fd._2892_ fd._3068_ fd._3112_ fd._3123_ VGND VGND VPWR VPWR fd._3134_ sky130_fd_sc_hd__a31o_1
XFILLER_226_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7147_ fd._2355_ fd._2360_ fd._2387_ fd._2388_ VGND VGND VPWR VPWR fd._2389_ sky130_fd_sc_hd__a31o_1
XFILLER_148_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_270_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_1606 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7078_ fd._2310_ fd._2312_ VGND VGND VPWR VPWR fd._2313_ sky130_fd_sc_hd__nor2_1
XFILLER_35_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_282_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6029_ fd._0972_ fd._1158_ VGND VGND VPWR VPWR fd._1159_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_254_1702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_274_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_249_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_259_1668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_project_wrapper_204 VGND VGND VPWR VPWR user_project_wrapper_204/HI la_data_out[82]
+ sky130_fd_sc_hd__conb_1
XFILLER_181_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_project_wrapper_215 VGND VGND VPWR VPWR user_project_wrapper_215/HI la_data_out[93]
+ sky130_fd_sc_hd__conb_1
XFILLER_103_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_project_wrapper_226 VGND VGND VPWR VPWR user_project_wrapper_226/HI la_data_out[104]
+ sky130_fd_sc_hd__conb_1
XFILLER_86_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_project_wrapper_237 VGND VGND VPWR VPWR user_project_wrapper_237/HI la_data_out[115]
+ sky130_fd_sc_hd__conb_1
Xuser_project_wrapper_248 VGND VGND VPWR VPWR user_project_wrapper_248/HI la_data_out[126]
+ sky130_fd_sc_hd__conb_1
XFILLER_5_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_project_wrapper_259 VGND VGND VPWR VPWR user_project_wrapper_259/HI wbs_dat_o[5]
+ sky130_fd_sc_hd__conb_1
XFILLER_190_1502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5400_ fd._0413_ fd._0466_ VGND VGND VPWR VPWR fd._0467_ sky130_fd_sc_hd__or2b_1
XFILLER_150_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6380_ fd._1371_ fd._1544_ VGND VGND VPWR VPWR fd._1545_ sky130_fd_sc_hd__xnor2_1
XTAP_6150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5331_ fd._0388_ fd._0390_ VGND VGND VPWR VPWR fd._0391_ sky130_fd_sc_hd__xnor2_1
XTAP_6183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_255_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5262_ fd._0113_ fd._0314_ VGND VGND VPWR VPWR fd._0315_ sky130_fd_sc_hd__xnor2_1
Xfd._8050_ fd._3364_ fd._3369_ fd._3375_ fd._3381_ VGND VGND VPWR VPWR fd._3382_ sky130_fd_sc_hd__and4_1
XFILLER_23_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4213_ fd._1451_ fd._1517_ VGND VGND VPWR VPWR fd._1528_ sky130_fd_sc_hd__nand2_1
XFILLER_188_1464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7001_ fd._2126_ fd._2222_ VGND VGND VPWR VPWR fd._2228_ sky130_fd_sc_hd__and2_1
XFILLER_149_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5193_ fd._0049_ fd._0237_ fd._0238_ VGND VGND VPWR VPWR fd._0239_ sky130_fd_sc_hd__o21ba_2
XFILLER_208_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4144_ fd._0758_ fd.a\[13\] VGND VGND VPWR VPWR fd._0769_ sky130_fd_sc_hd__nor2_1
XFILLER_51_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4075_ fd.b\[20\] fd._4071_ VGND VGND VPWR VPWR fd._0010_ sky130_fd_sc_hd__nor2_1
XFILLER_264_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_264_1396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7903_ fd._3047_ fd._3219_ fd._3077_ VGND VGND VPWR VPWR fd._3220_ sky130_fd_sc_hd__mux2_1
XFILLER_149_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7834_ fd._3141_ fd._3143_ VGND VGND VPWR VPWR fd._3144_ sky130_fd_sc_hd__xnor2_1
XFILLER_191_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7765_ fd._3066_ fd._3067_ VGND VGND VPWR VPWR fd._3069_ sky130_fd_sc_hd__or2b_1
XFILLER_117_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4977_ fd._3923_ fd._0001_ VGND VGND VPWR VPWR fd._0002_ sky130_fd_sc_hd__and2_1
XFILLER_118_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._6716_ fd._1842_ fd._1908_ fd._1911_ fd._1912_ fd._1914_ VGND VGND VPWR VPWR fd._1915_
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_156_1408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7696_ fd._2707_ fd._2798_ fd._2800_ VGND VGND VPWR VPWR fd._2993_ sky130_fd_sc_hd__a21oi_1
XFILLER_278_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6647_ fd._1699_ fd._1838_ fd._1813_ VGND VGND VPWR VPWR fd._1839_ sky130_fd_sc_hd__a21o_1
XFILLER_235_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6578_ fd._0437_ fd._1617_ VGND VGND VPWR VPWR fd._1763_ sky130_fd_sc_hd__and2_1
XFILLER_99_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5529_ fd._0469_ VGND VGND VPWR VPWR fd._0609_ sky130_fd_sc_hd__inv_2
XFILLER_41_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8248_ net75 net31 VGND VGND VPWR VPWR fd.b\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8179_ net77 fd.mc\[3\] VGND VGND VPWR VPWR fd.c\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_227_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_282_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout67 net69 VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_2
XFILLER_211_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_250_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_1547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_246_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4900_ fd._3688_ fd._3879_ fd._3880_ VGND VGND VPWR VPWR fd._3994_ sky130_fd_sc_hd__o21ai_1
XFILLER_35_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5880_ fd._0858_ VGND VGND VPWR VPWR fd._0995_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_173_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_259_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4831_ fd._3817_ fd._3924_ VGND VGND VPWR VPWR fd._3925_ sky130_fd_sc_hd__nand2_1
XFILLER_173_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7550_ fd._2645_ fd._2654_ VGND VGND VPWR VPWR fd._2832_ sky130_fd_sc_hd__nand2_1
XFILLER_138_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4762_ fd._3854_ fd._3855_ VGND VGND VPWR VPWR fd._3856_ sky130_fd_sc_hd__xnor2_1
XFILLER_170_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6501_ fd._1675_ fd._1677_ fd._1615_ VGND VGND VPWR VPWR fd._1678_ sky130_fd_sc_hd__o21ba_1
XFILLER_141_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7481_ fd._2377_ fd._2753_ fd._2754_ VGND VGND VPWR VPWR fd._2756_ sky130_fd_sc_hd__o21a_1
Xfd._4693_ fd._3786_ VGND VGND VPWR VPWR fd._3787_ sky130_fd_sc_hd__buf_8
XFILLER_142_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6432_ fd._1358_ fd._1601_ fd._1533_ VGND VGND VPWR VPWR fd._1602_ sky130_fd_sc_hd__mux2_1
XFILLER_116_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_269_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6363_ fd._1321_ fd._1423_ VGND VGND VPWR VPWR fd._1526_ sky130_fd_sc_hd__nand2_1
XFILLER_42_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8102_ fd._3420_ VGND VGND VPWR VPWR fd.mc\[18\] sky130_fd_sc_hd__clkbuf_1
Xfd._5314_ fd._0174_ fd._0371_ fd._0269_ VGND VGND VPWR VPWR fd._0372_ sky130_fd_sc_hd__mux2_1
XFILLER_83_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._6294_ fd._1177_ fd._1227_ fd._1174_ VGND VGND VPWR VPWR fd._1450_ sky130_fd_sc_hd__a21boi_1
XTAP_5290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8033_ fd._3086_ fd._3362_ fd._3241_ VGND VGND VPWR VPWR fd._3363_ sky130_fd_sc_hd__mux2_1
XFILLER_97_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_264_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5245_ fd._3708_ fd._0139_ VGND VGND VPWR VPWR fd._0297_ sky130_fd_sc_hd__and2_1
XFILLER_188_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5176_ fd._0220_ fd._0031_ fd._0067_ VGND VGND VPWR VPWR fd._0221_ sky130_fd_sc_hd__mux2_1
XFILLER_197_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4127_ fd.a\[10\] fd.b\[10\] VGND VGND VPWR VPWR fd._0582_ sky130_fd_sc_hd__and2b_1
XFILLER_240_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7817_ fd._2905_ fd._3125_ fd._3076_ VGND VGND VPWR VPWR fd._3126_ sky130_fd_sc_hd__mux2_1
XFILLER_69_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7748_ fd._3043_ fd._3048_ fd._3049_ VGND VGND VPWR VPWR fd._3050_ sky130_fd_sc_hd__and3_1
XFILLER_69_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_279_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7679_ fd._1722_ fd._2917_ VGND VGND VPWR VPWR fd._2974_ sky130_fd_sc_hd__nand2_1
XFILLER_121_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_230_ fd.c\[22\] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_1
XFILLER_23_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_1663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_284_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_250_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5030_ fd._0059_ VGND VGND VPWR VPWR fd._0060_ sky130_fd_sc_hd__buf_6
XFILLER_222_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_283_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._6981_ fd._2134_ fd._2140_ fd._2195_ fd._2204_ fd._2205_ VGND VGND VPWR VPWR fd._2206_
+ sky130_fd_sc_hd__o41a_1
XFILLER_92_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_261_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5932_ fd._2738_ fd._1051_ VGND VGND VPWR VPWR fd._1052_ sky130_fd_sc_hd__nand2_1
XFILLER_187_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5863_ fd._0885_ VGND VGND VPWR VPWR fd._0976_ sky130_fd_sc_hd__inv_2
XFILLER_31_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7602_ fd._2688_ fd._2809_ VGND VGND VPWR VPWR fd._2889_ sky130_fd_sc_hd__or2_1
Xfd._4814_ fd._3853_ fd._3899_ fd._3907_ fd._3904_ VGND VGND VPWR VPWR fd._3908_ sky130_fd_sc_hd__a31o_1
XFILLER_155_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5794_ fd._0898_ fd._0899_ VGND VGND VPWR VPWR fd._0900_ sky130_fd_sc_hd__and2_1
XFILLER_127_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7533_ fd._2677_ VGND VGND VPWR VPWR fd._2813_ sky130_fd_sc_hd__buf_6
XFILLER_5_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4745_ fd._3833_ fd._3838_ VGND VGND VPWR VPWR fd._3839_ sky130_fd_sc_hd__and2_1
XFILLER_192_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_272_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._7464_ fd._2735_ fd._2736_ VGND VGND VPWR VPWR fd._2737_ sky130_fd_sc_hd__and2_1
Xfd._4676_ fd._3617_ fd._3769_ VGND VGND VPWR VPWR fd._3770_ sky130_fd_sc_hd__nor2_1
XFILLER_269_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_256_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6415_ fd._0437_ fd._1423_ VGND VGND VPWR VPWR fd._1584_ sky130_fd_sc_hd__nand2_1
XFILLER_68_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7395_ fd._2494_ fd._2660_ fd._2499_ VGND VGND VPWR VPWR fd._2662_ sky130_fd_sc_hd__o21a_1
XFILLER_29_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_284_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_272_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6346_ fd._1303_ fd._1307_ fd._1339_ VGND VGND VPWR VPWR fd._1508_ sky130_fd_sc_hd__o21a_1
XFILLER_84_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput2 io_in[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_2
XFILLER_216_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_256_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_272_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6277_ fd._1296_ fd._1295_ fd._1422_ VGND VGND VPWR VPWR fd._1432_ sky130_fd_sc_hd__nand3b_1
XFILLER_37_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8016_ fd._1656_ fd._3126_ VGND VGND VPWR VPWR fd._3345_ sky130_fd_sc_hd__or2_1
XFILLER_77_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5228_ fd._2738_ fd._0276_ VGND VGND VPWR VPWR fd._0278_ sky130_fd_sc_hd__or2_1
XFILLER_225_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_244_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._5159_ fd._3972_ VGND VGND VPWR VPWR fd._0202_ sky130_fd_sc_hd__inv_2
XFILLER_240_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_279_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_8107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_251_1546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_259_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_1519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_230_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_213_ fd.c\[5\] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_1
XFILLER_169_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4530_ fd._3600_ fd._3606_ fd._3618_ fd._3623_ VGND VGND VPWR VPWR fd._3624_ sky130_fd_sc_hd__a31o_4
XFILLER_140_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4461_ fd._3553_ fd._3554_ fd.b\[11\] VGND VGND VPWR VPWR fd._3555_ sky130_fd_sc_hd__a21o_1
XFILLER_152_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6200_ fd._1322_ fd._1335_ fd._1346_ VGND VGND VPWR VPWR fd._1347_ sky130_fd_sc_hd__or3_1
XFILLER_254_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7180_ fd._2424_ VGND VGND VPWR VPWR fd._2425_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_66_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4392_ fd.b\[9\] VGND VGND VPWR VPWR fd._3469_ sky130_fd_sc_hd__buf_6
XFILLER_65_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6131_ fd._1268_ fd._1270_ VGND VGND VPWR VPWR fd._1271_ sky130_fd_sc_hd__xnor2_1
XFILLER_47_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6062_ fd._1190_ fd._1194_ fd._1169_ VGND VGND VPWR VPWR fd._1195_ sky130_fd_sc_hd__mux2_1
XFILLER_185_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_280_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_262_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5013_ fd._0039_ fd._0040_ VGND VGND VPWR VPWR fd._0041_ sky130_fd_sc_hd__nand2_1
XFILLER_179_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6964_ fd._1976_ fd._2185_ fd._2186_ fd._1585_ VGND VGND VPWR VPWR fd._2187_ sky130_fd_sc_hd__a211o_1
XFILLER_159_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._5915_ fd._1003_ fd._1007_ fd._1032_ VGND VGND VPWR VPWR fd._1034_ sky130_fd_sc_hd__or3_1
XFILLER_119_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._6895_ fd._2047_ VGND VGND VPWR VPWR fd._2112_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_175_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5846_ fd._0957_ VGND VGND VPWR VPWR fd._0958_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_116_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5777_ fd._0749_ fd._0881_ VGND VGND VPWR VPWR fd._0882_ sky130_fd_sc_hd__nand2_1
XFILLER_118_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7516_ fd._1872_ fd._2706_ VGND VGND VPWR VPWR fd._2795_ sky130_fd_sc_hd__nand2_1
Xfd._4728_ fd._1297_ fd._3820_ VGND VGND VPWR VPWR fd._3822_ sky130_fd_sc_hd__or2_1
XFILLER_143_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7447_ fd._2522_ VGND VGND VPWR VPWR fd._2719_ sky130_fd_sc_hd__clkinv_2
Xfd._4659_ fd._3581_ fd._3578_ fd._3579_ VGND VGND VPWR VPWR fd._3753_ sky130_fd_sc_hd__a21bo_1
XFILLER_130_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_257_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7378_ fd._2454_ fd._2642_ fd._2506_ VGND VGND VPWR VPWR fd._2643_ sky130_fd_sc_hd__and3_1
XFILLER_116_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_272_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6329_ fd._0965_ fd._1443_ VGND VGND VPWR VPWR fd._1489_ sky130_fd_sc_hd__or2_1
XFILLER_256_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_1596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_1615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_271_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_1659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_244_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_279_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_279_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_273_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_250_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_280_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_284_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_280_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_1461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5700_ fd._0477_ fd._0783_ fd._0460_ VGND VGND VPWR VPWR fd._0797_ sky130_fd_sc_hd__a21bo_1
XFILLER_156_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6680_ fd._1650_ fd._1873_ VGND VGND VPWR VPWR fd._1875_ sky130_fd_sc_hd__or2_1
XTAP_9150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5631_ fd._0708_ fd._0715_ fd._0719_ fd._0720_ VGND VGND VPWR VPWR fd._0721_ sky130_fd_sc_hd__o211ai_1
XFILLER_125_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5562_ fd._3883_ fd._0616_ VGND VGND VPWR VPWR fd._0645_ sky130_fd_sc_hd__nor2_1
XFILLER_98_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7301_ fd._0318_ fd._2550_ fd._2556_ fd._0821_ fd._2557_ VGND VGND VPWR VPWR fd._2558_
+ sky130_fd_sc_hd__a221o_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4513_ fd._2892_ fd._3068_ VGND VGND VPWR VPWR fd._3607_ sky130_fd_sc_hd__nand2_1
XTAP_7781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_285_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5493_ fd._0564_ fd._0568_ VGND VGND VPWR VPWR fd._0569_ sky130_fd_sc_hd__or2_1
XFILLER_152_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7232_ fd._2294_ VGND VGND VPWR VPWR fd._2482_ sky130_fd_sc_hd__clkinv_2
XFILLER_79_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4444_ fd._3536_ fd._3200_ fd._3537_ VGND VGND VPWR VPWR fd._3538_ sky130_fd_sc_hd__o21a_1
XFILLER_113_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7163_ fd._2220_ fd._2219_ VGND VGND VPWR VPWR fd._2406_ sky130_fd_sc_hd__or2b_1
XFILLER_113_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4375_ fd._1429_ fd._3299_ fd._3211_ VGND VGND VPWR VPWR fd._3310_ sky130_fd_sc_hd__mux2_2
XFILLER_238_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6114_ fd._1250_ fd._1251_ fd._1087_ VGND VGND VPWR VPWR fd._1252_ sky130_fd_sc_hd__a21oi_1
XFILLER_4_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7094_ fd._2329_ fd._2204_ VGND VGND VPWR VPWR fd._2330_ sky130_fd_sc_hd__xnor2_1
XFILLER_39_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_263_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6045_ fd._1174_ fd._1175_ VGND VGND VPWR VPWR fd._1177_ sky130_fd_sc_hd__and2_1
XFILLER_39_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7996_ fd._3149_ fd._3152_ fd._3177_ fd._3147_ VGND VGND VPWR VPWR fd._3323_ sky130_fd_sc_hd__o31ai_1
XFILLER_21_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6947_ fd._1585_ fd._1980_ VGND VGND VPWR VPWR fd._2169_ sky130_fd_sc_hd__nor2_1
XFILLER_174_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6878_ fd._1118_ VGND VGND VPWR VPWR fd._2093_ sky130_fd_sc_hd__buf_6
XFILLER_159_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5829_ fd._3905_ fd._0938_ VGND VGND VPWR VPWR fd._0939_ sky130_fd_sc_hd__nor2_1
XFILLER_143_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_270_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_249_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_244_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_281_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_267_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_1610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4160_ fd._0670_ fd._0692_ fd._0659_ VGND VGND VPWR VPWR fd._0945_ sky130_fd_sc_hd__a21oi_1
XFILLER_188_1679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_1643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_223_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4091_ fd.b\[6\] fd.a\[6\] VGND VGND VPWR VPWR fd._0186_ sky130_fd_sc_hd__xor2_1
XFILLER_50_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7850_ fd._2956_ fd._3161_ fd._3075_ VGND VGND VPWR VPWR fd._3162_ sky130_fd_sc_hd__mux2_1
XPHY_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6801_ fd._1793_ fd._1969_ VGND VGND VPWR VPWR fd._2008_ sky130_fd_sc_hd__nand2_1
XFILLER_12_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7781_ fd._3085_ VGND VGND VPWR VPWR fd._3086_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_121_1527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._4993_ fd._0017_ fd._0018_ VGND VGND VPWR VPWR fd._0019_ sky130_fd_sc_hd__xnor2_1
XFILLER_156_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6732_ fd._1600_ fd._1923_ VGND VGND VPWR VPWR fd._1932_ sky130_fd_sc_hd__and2_1
XFILLER_157_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6663_ fd._1680_ fd._1855_ fd._1720_ VGND VGND VPWR VPWR fd._1856_ sky130_fd_sc_hd__mux2_1
XFILLER_193_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_1461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_256_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5614_ fd._0501_ fd._0690_ fd._0532_ VGND VGND VPWR VPWR fd._0702_ sky130_fd_sc_hd__and3_1
XFILLER_154_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6594_ fd._1543_ fd._1779_ VGND VGND VPWR VPWR fd._1780_ sky130_fd_sc_hd__xnor2_1
XTAP_8290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5545_ fd._0625_ fd._0443_ VGND VGND VPWR VPWR fd._0627_ sky130_fd_sc_hd__and2b_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8264_ net67 net17 VGND VGND VPWR VPWR fd.b\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_234_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_269_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5476_ fd._0360_ fd._0356_ VGND VGND VPWR VPWR fd._0551_ sky130_fd_sc_hd__and2b_1
XFILLER_239_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7215_ fd._2454_ fd._2459_ fd._2462_ VGND VGND VPWR VPWR fd._2464_ sky130_fd_sc_hd__a21o_1
XFILLER_67_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4427_ fd._0219_ fd._3519_ VGND VGND VPWR VPWR fd._3521_ sky130_fd_sc_hd__nand2_1
Xfd._8195_ net75 fd.mc\[19\] VGND VGND VPWR VPWR fd.c\[19\] sky130_fd_sc_hd__dfxtp_2
XFILLER_82_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7146_ fd._0504_ fd._2354_ VGND VGND VPWR VPWR fd._2388_ sky130_fd_sc_hd__nor2_1
XFILLER_270_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4358_ fd.b\[21\] fd._3101_ VGND VGND VPWR VPWR fd._3123_ sky130_fd_sc_hd__and2_1
XFILLER_214_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_281_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7077_ fd._1507_ fd._2311_ VGND VGND VPWR VPWR fd._2312_ sky130_fd_sc_hd__nor2_1
XFILLER_74_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4289_ fd._1451_ fd._1517_ VGND VGND VPWR VPWR fd._2364_ sky130_fd_sc_hd__xnor2_1
XFILLER_263_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6028_ fd._0970_ fd._1157_ fd._1047_ VGND VGND VPWR VPWR fd._1158_ sky130_fd_sc_hd__and3b_1
XFILLER_62_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_282_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_263_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7979_ fd._2135_ fd._3302_ fd._3297_ fd._0504_ VGND VGND VPWR VPWR fd._3304_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_191_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_274_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_270_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_252_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_252_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_260_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_281_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_259_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_project_wrapper_205 VGND VGND VPWR VPWR user_project_wrapper_205/HI la_data_out[83]
+ sky130_fd_sc_hd__conb_1
XFILLER_177_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xuser_project_wrapper_216 VGND VGND VPWR VPWR user_project_wrapper_216/HI la_data_out[94]
+ sky130_fd_sc_hd__conb_1
XFILLER_120_1560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_227 VGND VGND VPWR VPWR user_project_wrapper_227/HI la_data_out[105]
+ sky130_fd_sc_hd__conb_1
XFILLER_138_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_project_wrapper_238 VGND VGND VPWR VPWR user_project_wrapper_238/HI la_data_out[116]
+ sky130_fd_sc_hd__conb_1
Xuser_project_wrapper_249 VGND VGND VPWR VPWR user_project_wrapper_249/HI la_data_out[127]
+ sky130_fd_sc_hd__conb_1
XFILLER_68_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_268_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_268_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5330_ fd._0074_ fd._0389_ VGND VGND VPWR VPWR fd._0390_ sky130_fd_sc_hd__nand2_1
XTAP_6173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5261_ fd._0119_ fd._0132_ VGND VGND VPWR VPWR fd._0314_ sky130_fd_sc_hd__nor2_1
XFILLER_188_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7000_ fd._2126_ fd._2222_ fd._2226_ fd._2124_ VGND VGND VPWR VPWR fd._2227_ sky130_fd_sc_hd__a211o_1
XTAP_4771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4212_ fd.a\[11\] fd._1506_ fd._1220_ VGND VGND VPWR VPWR fd._1517_ sky130_fd_sc_hd__mux2_1
XFILLER_97_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_252_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5192_ fd._0046_ fd._0237_ VGND VGND VPWR VPWR fd._0238_ sky130_fd_sc_hd__xnor2_1
XFILLER_184_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_1427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4143_ fd.b\[13\] VGND VGND VPWR VPWR fd._0758_ sky130_fd_sc_hd__inv_2
XFILLER_223_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4074_ fd.a\[20\] VGND VGND VPWR VPWR fd._4071_ sky130_fd_sc_hd__inv_2
XFILLER_260_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7902_ fd._3216_ fd._3218_ VGND VGND VPWR VPWR fd._3219_ sky130_fd_sc_hd__xor2_1
XFILLER_242_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7833_ fd._2934_ fd._3142_ VGND VGND VPWR VPWR fd._3143_ sky130_fd_sc_hd__nand2_1
XFILLER_121_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7764_ fd._2481_ fd._3065_ VGND VGND VPWR VPWR fd._3067_ sky130_fd_sc_hd__or2_1
Xfd._4976_ fd._3828_ fd._3922_ fd._3823_ VGND VGND VPWR VPWR fd._0001_ sky130_fd_sc_hd__o21ai_1
XFILLER_238_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_1436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6715_ fd._1833_ VGND VGND VPWR VPWR fd._1914_ sky130_fd_sc_hd__inv_2
XFILLER_219_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7695_ fd._2896_ fd._2989_ fd._2990_ VGND VGND VPWR VPWR fd._2992_ sky130_fd_sc_hd__a21oi_1
XFILLER_172_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6646_ fd._1431_ fd._1837_ VGND VGND VPWR VPWR fd._1838_ sky130_fd_sc_hd__xnor2_1
XFILLER_275_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6577_ fd._1015_ fd._1761_ VGND VGND VPWR VPWR fd._1762_ sky130_fd_sc_hd__and2_1
XFILLER_59_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5528_ fd._0476_ fd._0607_ VGND VGND VPWR VPWR fd._0608_ sky130_fd_sc_hd__or2_1
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8247_ net75 net30 VGND VGND VPWR VPWR fd.b\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_251_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_255_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5459_ fd._0502_ fd._0496_ VGND VGND VPWR VPWR fd._0532_ sky130_fd_sc_hd__or2b_1
XFILLER_67_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8178_ net77 fd.mc\[2\] VGND VGND VPWR VPWR fd.c\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_242_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7129_ fd._1585_ fd._2186_ VGND VGND VPWR VPWR fd._2369_ sky130_fd_sc_hd__nor2_1
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_282_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout68 net69 VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_2
XFILLER_52_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_260_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1690 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4830_ fd._2584_ fd._3816_ VGND VGND VPWR VPWR fd._3924_ sky130_fd_sc_hd__or2_1
XFILLER_31_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4761_ fd._3674_ fd._3700_ VGND VGND VPWR VPWR fd._3855_ sky130_fd_sc_hd__and2b_1
XFILLER_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6500_ fd._4055_ fd._1676_ VGND VGND VPWR VPWR fd._1677_ sky130_fd_sc_hd__xnor2_1
XFILLER_126_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7480_ fd._2377_ fd._2753_ fd._2754_ VGND VGND VPWR VPWR fd._2755_ sky130_fd_sc_hd__nor3_1
XFILLER_141_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4692_ fd._3772_ fd._3783_ fd._3785_ VGND VGND VPWR VPWR fd._3786_ sky130_fd_sc_hd__and3_1
XFILLER_253_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_269_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6431_ fd._1361_ fd._1413_ VGND VGND VPWR VPWR fd._1601_ sky130_fd_sc_hd__xnor2_1
XFILLER_79_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_268_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6362_ fd._1520_ fd._1524_ VGND VGND VPWR VPWR fd._1525_ sky130_fd_sc_hd__and2b_1
XFILLER_81_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8101_ fd._0061_ fd._0270_ fd._3411_ VGND VGND VPWR VPWR fd._3420_ sky130_fd_sc_hd__mux2_1
XFILLER_205_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5313_ fd._0168_ fd._0370_ VGND VGND VPWR VPWR fd._0371_ sky130_fd_sc_hd__xnor2_1
XFILLER_42_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_284_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6293_ fd._1260_ VGND VGND VPWR VPWR fd._1449_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_114_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8032_ fd._3210_ fd._3361_ VGND VGND VPWR VPWR fd._3362_ sky130_fd_sc_hd__xor2_1
XFILLER_42_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5244_ fd._0086_ fd._0294_ fd._0269_ VGND VGND VPWR VPWR fd._0295_ sky130_fd_sc_hd__mux2_1
XFILLER_23_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_266_1448 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5175_ fd._0025_ fd._0035_ VGND VGND VPWR VPWR fd._0220_ sky130_fd_sc_hd__xnor2_1
XFILLER_221_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4126_ fd.b\[10\] fd.a\[10\] VGND VGND VPWR VPWR fd._0571_ sky130_fd_sc_hd__and2b_1
XFILLER_51_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._7816_ fd._2908_ fd._3124_ VGND VGND VPWR VPWR fd._3125_ sky130_fd_sc_hd__xor2_1
XFILLER_117_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4959_ fd._4047_ fd._4051_ fd._4053_ VGND VGND VPWR VPWR fd._4054_ sky130_fd_sc_hd__a21o_1
XFILLER_238_1528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7747_ fd._1507_ fd._3047_ VGND VGND VPWR VPWR fd._3049_ sky130_fd_sc_hd__nand2_1
XFILLER_238_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7678_ fd._1219_ fd._2970_ VGND VGND VPWR VPWR fd._2973_ sky130_fd_sc_hd__and2_1
XFILLER_271_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6629_ fd._1817_ fd._1818_ fd._1813_ VGND VGND VPWR VPWR fd._1819_ sky130_fd_sc_hd__mux2_1
XFILLER_8_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_262_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_1602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1635 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_1657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_265_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._6980_ fd._2202_ fd._2131_ fd._2201_ VGND VGND VPWR VPWR fd._2205_ sky130_fd_sc_hd__o21bai_1
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5931_ fd._1049_ fd._1050_ fd._1047_ VGND VGND VPWR VPWR fd._1051_ sky130_fd_sc_hd__mux2_1
XFILLER_147_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5862_ fd._0884_ fd._0974_ VGND VGND VPWR VPWR fd._0975_ sky130_fd_sc_hd__nor2_1
XFILLER_200_1627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4813_ fd._3904_ fd._3906_ VGND VGND VPWR VPWR fd._3907_ sky130_fd_sc_hd__nor2_1
Xfd._7601_ fd._2692_ fd._2807_ VGND VGND VPWR VPWR fd._2888_ sky130_fd_sc_hd__nand2_1
XFILLER_122_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._5793_ fd._0708_ fd._0715_ VGND VGND VPWR VPWR fd._0899_ sky130_fd_sc_hd__nand2_1
XFILLER_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7532_ fd._2646_ fd._2811_ VGND VGND VPWR VPWR fd._2812_ sky130_fd_sc_hd__xnor2_1
XFILLER_127_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4744_ fd._3837_ fd._3720_ fd._3787_ VGND VGND VPWR VPWR fd._3838_ sky130_fd_sc_hd__mux2_1
XFILLER_196_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_269_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7463_ fd._2141_ fd._2734_ VGND VGND VPWR VPWR fd._2736_ sky130_fd_sc_hd__or2_1
XFILLER_102_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4675_ fd._3611_ fd._3768_ VGND VGND VPWR VPWR fd._3769_ sky130_fd_sc_hd__nand2_1
XFILLER_142_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_272_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6414_ fd._1015_ fd._1581_ VGND VGND VPWR VPWR fd._1582_ sky130_fd_sc_hd__and2_1
XFILLER_269_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7394_ fd._2624_ fd._2489_ fd._2487_ VGND VGND VPWR VPWR fd._2660_ sky130_fd_sc_hd__a21o_1
XFILLER_9_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6345_ fd._0479_ VGND VGND VPWR VPWR fd._1507_ sky130_fd_sc_hd__buf_6
XFILLER_256_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput3 io_in[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_2
XFILLER_84_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6276_ fd._0594_ VGND VGND VPWR VPWR fd._1431_ sky130_fd_sc_hd__buf_6
XFILLER_42_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8015_ fd._3190_ fd._3195_ fd._3196_ VGND VGND VPWR VPWR fd._3344_ sky130_fd_sc_hd__a21o_1
XFILLER_37_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5227_ fd._2738_ fd._0276_ VGND VGND VPWR VPWR fd._0277_ sky130_fd_sc_hd__nand2_1
XFILLER_224_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5158_ fd._4070_ fd._0006_ fd._0004_ VGND VGND VPWR VPWR fd._0201_ sky130_fd_sc_hd__a21o_1
XFILLER_209_1641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4109_ fd.b\[1\] fd.a\[1\] VGND VGND VPWR VPWR fd._0384_ sky130_fd_sc_hd__and2b_1
XFILLER_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5089_ fd._3688_ VGND VGND VPWR VPWR fd._0125_ sky130_fd_sc_hd__buf_6
XFILLER_240_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_279_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_279_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_74 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_251_1558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_251_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_274_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_1610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_212_ fd.c\[4\] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_1
XFILLER_204_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._4460_ fd._3498_ fd._3549_ fd._3552_ fd._0857_ VGND VGND VPWR VPWR fd._3554_ sky130_fd_sc_hd__a31o_1
XTAP_7996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4391_ fd._3376_ fd._3422_ fd._3430_ fd._3439_ fd._3449_ VGND VGND VPWR VPWR fd._3459_
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_238_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6130_ fd._1269_ fd._1101_ VGND VGND VPWR VPWR fd._1270_ sky130_fd_sc_hd__nor2_1
XFILLER_24_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6061_ fd._1191_ fd._1193_ VGND VGND VPWR VPWR fd._1194_ sky130_fd_sc_hd__xor2_1
XFILLER_18_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_267_1576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_262_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._5012_ fd._3947_ fd._3962_ VGND VGND VPWR VPWR fd._0040_ sky130_fd_sc_hd__nand2_1
XFILLER_206_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6963_ fd._1970_ fd._2175_ fd._2176_ fd._2178_ VGND VGND VPWR VPWR fd._2186_ sky130_fd_sc_hd__and4_1
XFILLER_119_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5914_ fd._1014_ fd._1020_ fd._1029_ fd._1030_ fd._1031_ VGND VGND VPWR VPWR fd._1032_
+ sky130_fd_sc_hd__a311oi_2
XFILLER_31_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6894_ fd._2043_ fd._2037_ VGND VGND VPWR VPWR fd._2110_ sky130_fd_sc_hd__and2b_1
XFILLER_200_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5845_ fd._0721_ fd._0954_ fd._0848_ fd._0955_ VGND VGND VPWR VPWR fd._0957_ sky130_fd_sc_hd__a31o_1
XFILLER_174_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5776_ fd._0880_ fd._0746_ VGND VGND VPWR VPWR fd._0881_ sky130_fd_sc_hd__nand2_1
XFILLER_157_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4727_ fd._1297_ fd._3820_ VGND VGND VPWR VPWR fd._3821_ sky130_fd_sc_hd__nand2_1
Xfd._7515_ fd._2728_ fd._2786_ fd._2791_ fd._2792_ VGND VGND VPWR VPWR fd._2794_ sky130_fd_sc_hd__o31a_2
XFILLER_118_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_276_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4658_ fd._3633_ fd._3750_ fd._3751_ VGND VGND VPWR VPWR fd._3752_ sky130_fd_sc_hd__a21o_1
Xfd._7446_ fd._2566_ fd._2717_ VGND VGND VPWR VPWR fd._2718_ sky130_fd_sc_hd__or2_1
XFILLER_285_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7377_ fd._1494_ fd._2439_ fd._2453_ VGND VGND VPWR VPWR fd._2642_ sky130_fd_sc_hd__nand3_1
XFILLER_131_1529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4589_ fd.b\[2\] fd._3534_ VGND VGND VPWR VPWR fd._3683_ sky130_fd_sc_hd__nor2_1
XFILLER_29_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_986 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6328_ fd._1319_ fd._1487_ VGND VGND VPWR VPWR fd._1488_ sky130_fd_sc_hd__nand2_1
XFILLER_84_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6259_ fd._0928_ fd._1409_ VGND VGND VPWR VPWR fd._1412_ sky130_fd_sc_hd__or2_1
XFILLER_168_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_225_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_1641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_273_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_284_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_1435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5630_ fd._0712_ VGND VGND VPWR VPWR fd._0720_ sky130_fd_sc_hd__inv_2
XFILLER_197_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_1632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_9173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_259_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5561_ fd._3883_ fd._0616_ VGND VGND VPWR VPWR fd._0644_ sky130_fd_sc_hd__and2_1
XFILLER_140_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4512_ fd._3604_ fd._3605_ VGND VGND VPWR VPWR fd._3606_ sky130_fd_sc_hd__and2_1
XTAP_7771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7300_ fd._1764_ fd._2505_ fd._2555_ fd._0821_ fd._1211_ VGND VGND VPWR VPWR fd._2557_
+ sky130_fd_sc_hd__o221a_1
XFILLER_79_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5492_ fd._0366_ fd._0567_ fd._0452_ VGND VGND VPWR VPWR fd._0568_ sky130_fd_sc_hd__mux2_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7231_ fd._1632_ VGND VGND VPWR VPWR fd._2481_ sky130_fd_sc_hd__buf_4
XFILLER_87_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._4443_ fd.b\[1\] VGND VGND VPWR VPWR fd._3537_ sky130_fd_sc_hd__clkinv_4
XFILLER_39_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_282_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_269_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7162_ fd._2212_ fd._2213_ VGND VGND VPWR VPWR fd._2405_ sky130_fd_sc_hd__nand2_1
XFILLER_43_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4374_ fd._2408_ fd._3288_ VGND VGND VPWR VPWR fd._3299_ sky130_fd_sc_hd__or2_1
XFILLER_253_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6113_ fd._0526_ fd._0988_ fd._1095_ VGND VGND VPWR VPWR fd._1251_ sky130_fd_sc_hd__a21oi_1
XFILLER_187_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_254_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7093_ fd._2131_ fd._2328_ VGND VGND VPWR VPWR fd._2329_ sky130_fd_sc_hd__or2_1
XFILLER_19_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6044_ fd._1172_ fd._1170_ VGND VGND VPWR VPWR fd._1175_ sky130_fd_sc_hd__or2_1
XFILLER_165_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_245_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_280_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7995_ fd._3318_ fd._3319_ fd._3320_ VGND VGND VPWR VPWR fd._3322_ sky130_fd_sc_hd__or3b_1
XFILLER_124_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6946_ fd._1976_ fd._2167_ VGND VGND VPWR VPWR fd._2168_ sky130_fd_sc_hd__nand2_1
XFILLER_276_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6877_ fd._2083_ fd._2091_ VGND VGND VPWR VPWR fd._2092_ sky130_fd_sc_hd__nor2_1
XFILLER_102_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5828_ fd._0694_ fd._0937_ fd._0848_ VGND VGND VPWR VPWR fd._0938_ sky130_fd_sc_hd__mux2_1
XFILLER_137_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5759_ fd._0479_ fd._0860_ VGND VGND VPWR VPWR fd._0862_ sky130_fd_sc_hd__nor2_1
XFILLER_157_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_1620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_257_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7429_ fd._2600_ fd._2599_ VGND VGND VPWR VPWR fd._2699_ sky130_fd_sc_hd__or2b_1
XFILLER_131_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_273_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_281_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_279_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_283_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_264_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_251_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4090_ fd._0120_ fd._0142_ fd._0153_ fd._0164_ VGND VGND VPWR VPWR fd._0175_ sky130_fd_sc_hd__a31o_1
XFILLER_17_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_1688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._6800_ fd._1788_ fd._2006_ VGND VGND VPWR VPWR fd._2007_ sky130_fd_sc_hd__xnor2_1
Xfd._4992_ fd._3808_ fd._3929_ VGND VGND VPWR VPWR fd._0018_ sky130_fd_sc_hd__or2_1
XFILLER_223_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7780_ fd._2891_ fd._3084_ fd._3076_ VGND VGND VPWR VPWR fd._3085_ sky130_fd_sc_hd__mux2_1
XFILLER_12_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_258_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6731_ fd._1173_ fd._1930_ VGND VGND VPWR VPWR fd._1931_ sky130_fd_sc_hd__nand2_1
XFILLER_117_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6662_ fd._1674_ fd._1854_ VGND VGND VPWR VPWR fd._1855_ sky130_fd_sc_hd__xnor2_1
XFILLER_158_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5613_ fd._0501_ fd._0690_ fd._0532_ VGND VGND VPWR VPWR fd._0701_ sky130_fd_sc_hd__a21oi_1
XFILLER_158_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6593_ fd._1547_ fd._1599_ VGND VGND VPWR VPWR fd._1779_ sky130_fd_sc_hd__and2_1
XFILLER_256_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._5544_ fd._0125_ fd._0442_ VGND VGND VPWR VPWR fd._0625_ sky130_fd_sc_hd__nor2_1
XFILLER_154_1348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8263_ net67 net16 VGND VGND VPWR VPWR fd.b\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_234_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5475_ fd._0540_ fd._0547_ fd._0548_ VGND VGND VPWR VPWR fd._0550_ sky130_fd_sc_hd__o21bai_1
XFILLER_113_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_269_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4426_ fd._0219_ fd._3519_ VGND VGND VPWR VPWR fd._3520_ sky130_fd_sc_hd__or2_1
XFILLER_239_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7214_ fd._2461_ VGND VGND VPWR VPWR fd._2462_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_255_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8194_ net76 fd.mc\[18\] VGND VGND VPWR VPWR fd.c\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_254_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7145_ fd._2367_ fd._2374_ fd._2383_ fd._2384_ fd._2385_ VGND VGND VPWR VPWR fd._2387_
+ sky130_fd_sc_hd__a311o_1
XFILLER_113_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4357_ fd.b\[21\] fd._3101_ VGND VGND VPWR VPWR fd._3112_ sky130_fd_sc_hd__or2_1
XFILLER_255_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7076_ fd._2307_ VGND VGND VPWR VPWR fd._2311_ sky130_fd_sc_hd__inv_2
Xfd._4288_ fd._2331_ fd._2342_ fd._1627_ VGND VGND VPWR VPWR fd._2353_ sky130_fd_sc_hd__o21a_1
XFILLER_169_1591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_263_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6027_ fd._0098_ fd._0892_ fd._0969_ VGND VGND VPWR VPWR fd._1157_ sky130_fd_sc_hd__or3_1
XFILLER_179_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7978_ fd._2135_ fd._3302_ VGND VGND VPWR VPWR fd._3303_ sky130_fd_sc_hd__nor2_1
XFILLER_120_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6929_ fd._1948_ fd._2148_ fd._2115_ VGND VGND VPWR VPWR fd._2149_ sky130_fd_sc_hd__mux2_1
XFILLER_136_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_274_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_270_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_274_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_249_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_265_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_260_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_281_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_206 VGND VGND VPWR VPWR user_project_wrapper_206/HI la_data_out[84]
+ sky130_fd_sc_hd__conb_1
XFILLER_154_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_217 VGND VGND VPWR VPWR user_project_wrapper_217/HI la_data_out[95]
+ sky130_fd_sc_hd__conb_1
Xuser_project_wrapper_228 VGND VGND VPWR VPWR user_project_wrapper_228/HI la_data_out[106]
+ sky130_fd_sc_hd__conb_1
XFILLER_68_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_project_wrapper_239 VGND VGND VPWR VPWR user_project_wrapper_239/HI la_data_out[117]
+ sky130_fd_sc_hd__conb_1
XFILLER_153_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_253_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_270_1572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_283_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5260_ fd._0112_ VGND VGND VPWR VPWR fd._0313_ sky130_fd_sc_hd__clkinvlp_2
XTAP_5473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4211_ fd._0516_ fd._1495_ VGND VGND VPWR VPWR fd._1506_ sky130_fd_sc_hd__xnor2_1
XTAP_4761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5191_ fd._0038_ fd._0041_ fd._0039_ VGND VGND VPWR VPWR fd._0237_ sky130_fd_sc_hd__o21a_1
XTAP_4783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4142_ fd.b\[13\] fd._0736_ VGND VGND VPWR VPWR fd._0747_ sky130_fd_sc_hd__nor2_1
XFILLER_40_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_251_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4073_ fd.a\[22\] fd._4049_ VGND VGND VPWR VPWR fd._4060_ sky130_fd_sc_hd__or2_1
XFILLER_36_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_260_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_260_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7901_ fd._0768_ fd._3042_ fd._3217_ VGND VGND VPWR VPWR fd._3218_ sky130_fd_sc_hd__o21ba_1
XFILLER_149_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._7832_ fd._2533_ fd._2933_ VGND VGND VPWR VPWR fd._3142_ sky130_fd_sc_hd__or2_1
XFILLER_73_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7763_ fd._2481_ fd._3065_ VGND VGND VPWR VPWR fd._3066_ sky130_fd_sc_hd__and2_1
Xfd._4975_ fd._2584_ VGND VGND VPWR VPWR fd._0000_ sky130_fd_sc_hd__buf_6
XFILLER_172_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6714_ fd._1834_ fd._1824_ VGND VGND VPWR VPWR fd._1912_ sky130_fd_sc_hd__and2b_1
XFILLER_195_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7694_ fd._2093_ fd._2899_ fd._2988_ VGND VGND VPWR VPWR fd._2990_ sky130_fd_sc_hd__and3_1
XFILLER_132_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6645_ fd._1699_ fd._1702_ VGND VGND VPWR VPWR fd._1837_ sky130_fd_sc_hd__xor2_1
XFILLER_144_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6576_ fd._1588_ fd._1760_ fd._1719_ VGND VGND VPWR VPWR fd._1761_ sky130_fd_sc_hd__mux2_1
XFILLER_98_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5527_ fd._0026_ fd._0475_ VGND VGND VPWR VPWR fd._0607_ sky130_fd_sc_hd__and2_1
XFILLER_80_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8246_ net75 net29 VGND VGND VPWR VPWR fd.b\[6\] sky130_fd_sc_hd__dfxtp_2
XFILLER_41_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5458_ fd._0526_ fd._0530_ VGND VGND VPWR VPWR fd._0531_ sky130_fd_sc_hd__or2_1
XFILLER_80_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4409_ fd._1847_ fd._2023_ fd._2045_ VGND VGND VPWR VPWR fd._3503_ sky130_fd_sc_hd__a21oi_1
XFILLER_167_1506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5389_ fd._0454_ VGND VGND VPWR VPWR fd._0455_ sky130_fd_sc_hd__inv_2
XFILLER_167_1517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8177_ net77 fd.mc\[1\] VGND VGND VPWR VPWR fd.c\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_269_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_255_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7128_ fd._2179_ fd._2180_ fd._2183_ VGND VGND VPWR VPWR fd._2368_ sky130_fd_sc_hd__a21o_1
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_282_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7059_ fd._2066_ fd._2104_ VGND VGND VPWR VPWR fd._2292_ sky130_fd_sc_hd__nor2_1
XFILLER_126_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout69 net33 VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_6
XFILLER_22_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_276_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_276_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_276_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_1578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_259_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_1702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4760_ fd._3682_ fd._3699_ fd._3680_ VGND VGND VPWR VPWR fd._3854_ sky130_fd_sc_hd__o21ai_1
XFILLER_155_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4691_ fd._3628_ fd._3752_ fd._3756_ fd._3784_ fd._3782_ VGND VGND VPWR VPWR fd._3785_
+ sky130_fd_sc_hd__a2111o_1
XFILLER_177_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_272_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_253_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6430_ fd._0916_ VGND VGND VPWR VPWR fd._1600_ sky130_fd_sc_hd__buf_4
XFILLER_155_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6361_ fd._1522_ fd._1523_ VGND VGND VPWR VPWR fd._1524_ sky130_fd_sc_hd__and2_1
XFILLER_150_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_268_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8100_ fd._3419_ VGND VGND VPWR VPWR fd.mc\[17\] sky130_fd_sc_hd__clkbuf_1
XFILLER_49_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5312_ fd._0176_ fd._0173_ VGND VGND VPWR VPWR fd._0370_ sky130_fd_sc_hd__and2b_1
Xfd._6292_ fd._1445_ fd._1447_ fd._1422_ VGND VGND VPWR VPWR fd._1448_ sky130_fd_sc_hd__mux2_1
XTAP_5270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5243_ fd._0146_ fd._0293_ VGND VGND VPWR VPWR fd._0294_ sky130_fd_sc_hd__xnor2_1
Xfd._8031_ fd._3093_ fd._3096_ fd._3207_ fd._3208_ VGND VGND VPWR VPWR fd._3361_ sky130_fd_sc_hd__a31oi_1
XFILLER_252_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5174_ fd._0217_ VGND VGND VPWR VPWR fd._0218_ sky130_fd_sc_hd__clkinv_4
XFILLER_188_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4125_ fd._0527_ fd._0549_ VGND VGND VPWR VPWR fd._0560_ sky130_fd_sc_hd__nand2_1
XFILLER_166_1550 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_264_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_1545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_260_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7815_ fd._2920_ fd._2976_ VGND VGND VPWR VPWR fd._3124_ sky130_fd_sc_hd__nand2_1
XFILLER_118_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7746_ fd._1507_ fd._3047_ VGND VGND VPWR VPWR fd._3048_ sky130_fd_sc_hd__or2_1
XFILLER_121_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4958_ fd._0758_ fd._4052_ VGND VGND VPWR VPWR fd._4053_ sky130_fd_sc_hd__nor2_1
XFILLER_195_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_279_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._7677_ fd._2919_ fd._2912_ VGND VGND VPWR VPWR fd._2972_ sky130_fd_sc_hd__or2b_1
XFILLER_47_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4889_ fd._3874_ fd._3881_ VGND VGND VPWR VPWR fd._3983_ sky130_fd_sc_hd__and2_1
XFILLER_99_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6628_ fd._1806_ fd._1711_ VGND VGND VPWR VPWR fd._1818_ sky130_fd_sc_hd__xor2_1
XFILLER_86_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6559_ fd._1739_ fd._1741_ VGND VGND VPWR VPWR fd._1742_ sky130_fd_sc_hd__xnor2_1
XFILLER_59_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8229_ net70 net14 VGND VGND VPWR VPWR fd.a\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_255_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_270_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_273_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_261_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_261_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5930_ fd._1041_ fd._0982_ VGND VGND VPWR VPWR fd._1050_ sky130_fd_sc_hd__xnor2_1
XFILLER_187_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5861_ fd._0594_ fd._0883_ VGND VGND VPWR VPWR fd._0974_ sky130_fd_sc_hd__and2_1
XFILLER_139_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7600_ fd._2885_ fd._2886_ VGND VGND VPWR VPWR fd._2887_ sky130_fd_sc_hd__nand2_1
XFILLER_274_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4812_ fd._3905_ fd._3903_ VGND VGND VPWR VPWR fd._3906_ sky130_fd_sc_hd__nor2_1
XFILLER_31_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5792_ fd._0708_ fd._0715_ VGND VGND VPWR VPWR fd._0898_ sky130_fd_sc_hd__or2_1
XFILLER_154_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_259_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7531_ fd._2653_ fd._2652_ VGND VGND VPWR VPWR fd._2811_ sky130_fd_sc_hd__or2b_1
XFILLER_5_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4743_ fd._3834_ fd._3836_ VGND VGND VPWR VPWR fd._3837_ sky130_fd_sc_hd__xnor2_1
XFILLER_196_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7462_ fd._2141_ fd._2734_ VGND VGND VPWR VPWR fd._2735_ sky130_fd_sc_hd__nand2_1
Xfd._4674_ fd._3613_ fd._3761_ VGND VGND VPWR VPWR fd._3768_ sky130_fd_sc_hd__or2b_1
XFILLER_269_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6413_ fd._1576_ fd._1580_ fd._1533_ VGND VGND VPWR VPWR fd._1581_ sky130_fd_sc_hd__mux2_1
XFILLER_284_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7393_ fd._1507_ fd._2630_ fd._2636_ fd._2658_ VGND VGND VPWR VPWR fd._2659_ sky130_fd_sc_hd__a22o_1
XFILLER_110_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_284_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._6344_ fd._1425_ fd._1430_ fd._1503_ fd._1504_ fd._1088_ VGND VGND VPWR VPWR fd._1505_
+ sky130_fd_sc_hd__a32o_1
XFILLER_81_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput4 io_in[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_2
XFILLER_237_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6275_ fd._0131_ fd._1428_ VGND VGND VPWR VPWR fd._1430_ sky130_fd_sc_hd__or2_1
XFILLER_168_1612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8014_ fd._1330_ fd._3340_ VGND VGND VPWR VPWR fd._3342_ sky130_fd_sc_hd__and2_1
XFILLER_252_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5226_ fd._0222_ fd._0275_ fd._0270_ VGND VGND VPWR VPWR fd._0276_ sky130_fd_sc_hd__mux2_1
XFILLER_224_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5157_ fd._0075_ fd._0199_ VGND VGND VPWR VPWR fd._0200_ sky130_fd_sc_hd__or2_1
XFILLER_51_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4108_ fd.b\[1\] fd.a\[1\] VGND VGND VPWR VPWR fd._0373_ sky130_fd_sc_hd__xnor2_1
Xfd._5088_ fd._0050_ fd._0052_ fd._0057_ fd._0123_ VGND VGND VPWR VPWR fd._0124_ sky130_fd_sc_hd__a31oi_1
XFILLER_221_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_1686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7729_ fd._3028_ fd._2829_ fd._2849_ VGND VGND VPWR VPWR fd._3029_ sky130_fd_sc_hd__a21o_1
XFILLER_279_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_1662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_255_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_211_ fd.c\[3\] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_2
XFILLER_243_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_9300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_266_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4390_ fd.b\[14\] fd._3310_ VGND VGND VPWR VPWR fd._3449_ sky130_fd_sc_hd__xnor2_2
XFILLER_215_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_281_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6060_ fd._1020_ fd._1192_ VGND VGND VPWR VPWR fd._1193_ sky130_fd_sc_hd__and2_1
XFILLER_20_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5011_ fd._3947_ fd._3962_ VGND VGND VPWR VPWR fd._0039_ sky130_fd_sc_hd__or2_1
XFILLER_34_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_261_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6962_ fd._2175_ fd._2176_ fd._2178_ fd._2182_ VGND VGND VPWR VPWR fd._2185_ sky130_fd_sc_hd__a31o_1
XFILLER_147_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5913_ fd._0807_ fd._1005_ VGND VGND VPWR VPWR fd._1031_ sky130_fd_sc_hd__nor2_1
XFILLER_186_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6893_ fd._0768_ fd._2041_ VGND VGND VPWR VPWR fd._2109_ sky130_fd_sc_hd__xnor2_2
XFILLER_31_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_278_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_1602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5844_ fd._0660_ fd._0848_ VGND VGND VPWR VPWR fd._0955_ sky130_fd_sc_hd__nor2_1
XFILLER_116_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5775_ fd._0000_ fd._0744_ fd._0748_ VGND VGND VPWR VPWR fd._0880_ sky130_fd_sc_hd__a21o_1
XFILLER_142_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7514_ fd._2326_ fd._2790_ VGND VGND VPWR VPWR fd._2792_ sky130_fd_sc_hd__or2_1
Xfd._4726_ fd._3819_ fd._3736_ fd._3788_ VGND VGND VPWR VPWR fd._3820_ sky130_fd_sc_hd__mux2_1
XFILLER_192_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7445_ fd._2514_ fd._2715_ fd._2676_ VGND VGND VPWR VPWR fd._2717_ sky130_fd_sc_hd__mux2_1
XFILLER_285_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._4657_ fd.b\[19\] fd._3627_ VGND VGND VPWR VPWR fd._3751_ sky130_fd_sc_hd__and2_1
XFILLER_233_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7376_ fd._2465_ fd._2640_ VGND VGND VPWR VPWR fd._2641_ sky130_fd_sc_hd__or2_1
XFILLER_9_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4588_ fd._3680_ fd._3681_ VGND VGND VPWR VPWR fd._3682_ sky130_fd_sc_hd__nand2_1
XFILLER_111_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_285_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_250_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_284_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6327_ fd._1240_ fd._1486_ fd._1422_ VGND VGND VPWR VPWR fd._1487_ sky130_fd_sc_hd__mux2_1
XFILLER_256_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_272_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6258_ fd._1219_ fd._1410_ VGND VGND VPWR VPWR fd._1411_ sky130_fd_sc_hd__nor2_1
XFILLER_77_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_271_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5209_ fd._0253_ fd._0255_ fd._0256_ VGND VGND VPWR VPWR fd._0257_ sky130_fd_sc_hd__a21oi_1
XFILLER_198_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6189_ fd._1165_ fd._1332_ VGND VGND VPWR VPWR fd._1335_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_244_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1615 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_279_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_268_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_263_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_212_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_9130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_9174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_9196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5560_ fd._0623_ fd._0641_ fd._0642_ VGND VGND VPWR VPWR fd._0643_ sky130_fd_sc_hd__a21oi_1
XFILLER_139_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4511_ fd.b\[21\] fd._3603_ VGND VGND VPWR VPWR fd._3605_ sky130_fd_sc_hd__or2_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5491_ fd._0565_ fd._0566_ VGND VGND VPWR VPWR fd._0567_ sky130_fd_sc_hd__nor2_1
XFILLER_79_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7230_ fd._2472_ fd._2479_ VGND VGND VPWR VPWR fd._2480_ sky130_fd_sc_hd__or2b_1
XFILLER_267_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4442_ fd.b\[0\] VGND VGND VPWR VPWR fd._3536_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_6_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_266_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7161_ fd._2399_ fd._2403_ fd._1797_ fd._2402_ VGND VGND VPWR VPWR fd._2404_ sky130_fd_sc_hd__o2bb2a_1
Xfd._4373_ fd._1528_ fd._2375_ fd._2397_ VGND VGND VPWR VPWR fd._3288_ sky130_fd_sc_hd__and3_1
XFILLER_238_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_254_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6112_ fd._1092_ VGND VGND VPWR VPWR fd._1250_ sky130_fd_sc_hd__inv_2
XFILLER_282_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7092_ fd._2134_ fd._2140_ fd._2195_ VGND VGND VPWR VPWR fd._2328_ sky130_fd_sc_hd__nor3_1
XFILLER_207_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_267_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_253_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6043_ fd._1173_ fd._1170_ VGND VGND VPWR VPWR fd._1174_ sky130_fd_sc_hd__nand2_1
XFILLER_165_1615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7994_ fd._1797_ fd._3313_ VGND VGND VPWR VPWR fd._3320_ sky130_fd_sc_hd__nand2_1
XFILLER_148_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._6945_ fd._1969_ fd._1971_ fd._1974_ VGND VGND VPWR VPWR fd._2167_ sky130_fd_sc_hd__a21o_1
XFILLER_174_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6876_ fd._1645_ fd._2090_ VGND VGND VPWR VPWR fd._2091_ sky130_fd_sc_hd__nor2_1
XFILLER_159_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5827_ fd._0936_ fd._0698_ VGND VGND VPWR VPWR fd._0937_ sky130_fd_sc_hd__xnor2_1
XFILLER_157_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5758_ fd._0479_ fd._0860_ VGND VGND VPWR VPWR fd._0861_ sky130_fd_sc_hd__nand2_1
XFILLER_103_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4709_ fd._1352_ fd._3802_ VGND VGND VPWR VPWR fd._3803_ sky130_fd_sc_hd__or2_1
XFILLER_118_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5689_ fd._0459_ fd._0784_ fd._0651_ VGND VGND VPWR VPWR fd._0785_ sky130_fd_sc_hd__mux2_1
XFILLER_272_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_1676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7428_ fd._1645_ fd._2697_ VGND VGND VPWR VPWR fd._2698_ sky130_fd_sc_hd__nand2_1
XFILLER_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_270_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_268_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7359_ fd._2616_ fd._2621_ VGND VGND VPWR VPWR fd._2622_ sky130_fd_sc_hd__xnor2_1
XFILLER_29_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_268_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_272_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_272_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_279_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_253_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_251_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_264_1514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_251_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_1678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4991_ fd._3813_ fd._3928_ VGND VGND VPWR VPWR fd._0017_ sky130_fd_sc_hd__nor2_1
XFILLER_156_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6730_ fd._1735_ fd._1929_ fd._1917_ VGND VGND VPWR VPWR fd._1930_ sky130_fd_sc_hd__mux2_1
XFILLER_156_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6661_ fd._1683_ fd._1681_ VGND VGND VPWR VPWR fd._1854_ sky130_fd_sc_hd__nor2_1
XFILLER_172_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5612_ fd._0669_ fd._0676_ fd._0688_ fd._0698_ fd._0699_ VGND VGND VPWR VPWR fd._0700_
+ sky130_fd_sc_hd__a41o_1
XTAP_8270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._6592_ fd._1746_ fd._1750_ fd._1776_ fd._1777_ fd._1744_ VGND VGND VPWR VPWR fd._1778_
+ sky130_fd_sc_hd__o311a_1
XFILLER_119_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5543_ fd._4011_ fd._0444_ VGND VGND VPWR VPWR fd._0624_ sky130_fd_sc_hd__nor2_1
XFILLER_234_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._8262_ net76 net15 VGND VGND VPWR VPWR fd.b\[22\] sky130_fd_sc_hd__dfxtp_2
XFILLER_234_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5474_ fd._3716_ fd._0546_ VGND VGND VPWR VPWR fd._0548_ sky130_fd_sc_hd__and2_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7213_ fd._2434_ fd._2460_ VGND VGND VPWR VPWR fd._2461_ sky130_fd_sc_hd__and2_1
XFILLER_269_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4425_ fd._1880_ fd._3518_ fd._3200_ VGND VGND VPWR VPWR fd._3519_ sky130_fd_sc_hd__mux2_1
XFILLER_66_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8193_ net76 fd.mc\[17\] VGND VGND VPWR VPWR fd.c\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_230_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_212_1671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7144_ fd._1559_ fd._2359_ VGND VGND VPWR VPWR fd._2385_ sky130_fd_sc_hd__nor2_1
XFILLER_66_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4356_ fd._4071_ fd._3090_ fd._1231_ VGND VGND VPWR VPWR fd._3101_ sky130_fd_sc_hd__mux2_1
XFILLER_82_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_270_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7075_ fd._2308_ VGND VGND VPWR VPWR fd._2310_ sky130_fd_sc_hd__inv_2
XFILLER_35_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4287_ fd._0857_ fd._1605_ VGND VGND VPWR VPWR fd._2342_ sky130_fd_sc_hd__xnor2_2
XFILLER_208_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6026_ fd._1148_ fd._1153_ fd._1155_ VGND VGND VPWR VPWR fd._1156_ sky130_fd_sc_hd__a21o_1
XFILLER_78_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_280_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._7977_ fd._3146_ fd._3301_ fd._3239_ VGND VGND VPWR VPWR fd._3302_ sky130_fd_sc_hd__mux2_1
XFILLER_72_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6928_ fd._2146_ fd._2147_ VGND VGND VPWR VPWR fd._2148_ sky130_fd_sc_hd__xor2_1
XFILLER_11_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_276_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6859_ fd._1894_ fd._2071_ fd._1917_ VGND VGND VPWR VPWR fd._2072_ sky130_fd_sc_hd__mux2_1
XFILLER_151_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_249_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_281_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_281_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_207 VGND VGND VPWR VPWR user_project_wrapper_207/HI la_data_out[85]
+ sky130_fd_sc_hd__conb_1
XFILLER_193_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_218 VGND VGND VPWR VPWR user_project_wrapper_218/HI la_data_out[96]
+ sky130_fd_sc_hd__conb_1
XFILLER_257_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_229 VGND VGND VPWR VPWR user_project_wrapper_229/HI la_data_out[107]
+ sky130_fd_sc_hd__conb_1
XFILLER_68_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_283_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4210_ fd._0593_ fd._1484_ fd._0571_ VGND VGND VPWR VPWR fd._1495_ sky130_fd_sc_hd__a21o_1
XFILLER_236_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5190_ fd._0067_ fd._0121_ fd._0124_ VGND VGND VPWR VPWR fd._0236_ sky130_fd_sc_hd__a21o_1
XFILLER_149_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._4141_ fd.a\[13\] VGND VGND VPWR VPWR fd._0736_ sky130_fd_sc_hd__inv_2
XFILLER_252_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4072_ fd.b\[22\] VGND VGND VPWR VPWR fd._4049_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_210_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_260_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7900_ fd._3043_ fd._3074_ VGND VGND VPWR VPWR fd._3217_ sky130_fd_sc_hd__and2_1
XFILLER_17_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_1631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_242_1664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._7831_ fd._2943_ fd._2962_ fd._2963_ VGND VGND VPWR VPWR fd._3141_ sky130_fd_sc_hd__a21o_1
XFILLER_242_1675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_277_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7762_ fd._2879_ fd._3062_ fd._3064_ VGND VGND VPWR VPWR fd._3065_ sky130_fd_sc_hd__a21oi_1
XFILLER_117_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4974_ fd._4062_ fd._4068_ fd._4069_ VGND VGND VPWR VPWR fd._4070_ sky130_fd_sc_hd__a21boi_2
XFILLER_12_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6713_ fd._1909_ fd._1910_ VGND VGND VPWR VPWR fd._1911_ sky130_fd_sc_hd__nor2_1
XFILLER_117_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7693_ fd._2899_ fd._2988_ fd._2093_ VGND VGND VPWR VPWR fd._2989_ sky130_fd_sc_hd__a21o_1
XFILLER_12_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6644_ fd._1824_ fd._1829_ fd._1833_ fd._1834_ VGND VGND VPWR VPWR fd._1835_ sky130_fd_sc_hd__a211o_2
XFILLER_28_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6575_ fd._1590_ fd._1758_ VGND VGND VPWR VPWR fd._1760_ sky130_fd_sc_hd__xnor2_1
XFILLER_141_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_259_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5526_ fd._0482_ fd._0600_ fd._0605_ VGND VGND VPWR VPWR fd._0606_ sky130_fd_sc_hd__a21oi_2
XFILLER_141_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_246_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8245_ net72 net28 VGND VGND VPWR VPWR fd.b\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_239_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_255_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_251_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5457_ fd._0308_ fd._0529_ fd._0452_ VGND VGND VPWR VPWR fd._0530_ sky130_fd_sc_hd__mux2_1
XFILLER_171_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._4408_ fd._1682_ fd._3501_ fd._3200_ VGND VGND VPWR VPWR fd._3502_ sky130_fd_sc_hd__mux2_1
XFILLER_228_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8176_ net77 fd.mc\[0\] VGND VGND VPWR VPWR fd.c\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5388_ fd._0276_ fd._0451_ fd._0453_ VGND VGND VPWR VPWR fd._0454_ sky130_fd_sc_hd__mux2_2
XFILLER_270_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_265_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7127_ fd._1751_ fd._2366_ VGND VGND VPWR VPWR fd._2367_ sky130_fd_sc_hd__nand2_1
Xfd._4339_ fd._1033_ fd._2903_ fd._1220_ VGND VGND VPWR VPWR fd._2914_ sky130_fd_sc_hd__mux2_1
XFILLER_208_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_1504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7058_ fd._2258_ fd._2261_ fd._2290_ fd._2256_ VGND VGND VPWR VPWR fd._2291_ sky130_fd_sc_hd__a31o_1
XFILLER_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6009_ fd._0894_ fd._1136_ fd._1046_ VGND VGND VPWR VPWR fd._1137_ sky130_fd_sc_hd__mux2_1
XFILLER_195_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_278_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_265_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_1506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_1517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4690_ fd._3777_ fd._3778_ VGND VGND VPWR VPWR fd._3784_ sky130_fd_sc_hd__or2b_1
XFILLER_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_284_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6360_ fd._0786_ fd._1521_ VGND VGND VPWR VPWR fd._1523_ sky130_fd_sc_hd__nand2_1
XFILLER_123_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5311_ fd._0292_ fd._0361_ fd._0368_ fd._0365_ VGND VGND VPWR VPWR fd._0369_ sky130_fd_sc_hd__a31o_1
XFILLER_237_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_283_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6291_ fd._1267_ fd._1446_ VGND VGND VPWR VPWR fd._1447_ sky130_fd_sc_hd__xnor2_1
XTAP_5260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._8030_ fd._3357_ fd._3342_ fd._3355_ fd._3359_ VGND VGND VPWR VPWR fd._3360_ sky130_fd_sc_hd__o22ai_1
XFILLER_7_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5242_ fd._0136_ fd._0140_ fd._0144_ VGND VGND VPWR VPWR fd._0293_ sky130_fd_sc_hd__o21ai_1
XTAP_5293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5173_ fd._0215_ fd._0216_ VGND VGND VPWR VPWR fd._0217_ sky130_fd_sc_hd__or2_1
XFILLER_184_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_251_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4124_ fd.b\[9\] fd._0538_ VGND VGND VPWR VPWR fd._0549_ sky130_fd_sc_hd__nand2_1
XFILLER_264_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_264_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_260_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_277_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7814_ fd._3110_ fd._3117_ fd._3121_ VGND VGND VPWR VPWR fd._3122_ sky130_fd_sc_hd__or3_1
XFILLER_118_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7745_ fd._3044_ fd._3045_ fd._2877_ VGND VGND VPWR VPWR fd._3047_ sky130_fd_sc_hd__mux2_1
Xfd._4957_ fd._4050_ VGND VGND VPWR VPWR fd._4052_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_118_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7676_ fd._1219_ fd._2970_ VGND VGND VPWR VPWR fd._2971_ sky130_fd_sc_hd__or2_1
XFILLER_278_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4888_ fd._3469_ fd._3975_ fd._3981_ VGND VGND VPWR VPWR fd._3982_ sky130_fd_sc_hd__a21o_1
XFILLER_275_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6627_ fd._1630_ VGND VGND VPWR VPWR fd._1817_ sky130_fd_sc_hd__clkinv_2
XFILLER_138_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6558_ fd._1740_ fd._1595_ VGND VGND VPWR VPWR fd._1741_ sky130_fd_sc_hd__nor2_1
XFILLER_134_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_247_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5509_ fd._0381_ fd._0586_ VGND VGND VPWR VPWR fd._0587_ sky130_fd_sc_hd__xnor2_1
XFILLER_262_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6489_ fd._0758_ fd._1664_ VGND VGND VPWR VPWR fd._1665_ sky130_fd_sc_hd__nand2_1
XFILLER_132_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8228_ net70 net13 VGND VGND VPWR VPWR fd.a\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_216_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_255_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8159_ fd._3466_ fd._3472_ VGND VGND VPWR VPWR fd._3474_ sky130_fd_sc_hd__and2_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_282_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_243_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_265_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5860_ fd._0098_ fd._0892_ fd._0969_ fd._0972_ VGND VGND VPWR VPWR fd._0973_ sky130_fd_sc_hd__o31a_1
XFILLER_128_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4811_ fd._0857_ VGND VGND VPWR VPWR fd._3905_ sky130_fd_sc_hd__buf_6
XFILLER_139_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5791_ fd._0895_ fd._0896_ VGND VGND VPWR VPWR fd._0897_ sky130_fd_sc_hd__nor2_1
XFILLER_170_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7530_ fd._2692_ fd._2807_ fd._2809_ VGND VGND VPWR VPWR fd._2810_ sky130_fd_sc_hd__a21oi_1
Xfd._4742_ fd._3835_ fd._3721_ VGND VGND VPWR VPWR fd._3836_ sky130_fd_sc_hd__nor2_1
XFILLER_155_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_272_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7461_ fd._2729_ fd._2733_ fd._2676_ VGND VGND VPWR VPWR fd._2734_ sky130_fd_sc_hd__mux2_1
Xfd._4673_ fd.b\[22\] fd._3766_ VGND VGND VPWR VPWR fd._3767_ sky130_fd_sc_hd__nor2_1
XFILLER_142_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6412_ fd._1577_ fd._1579_ VGND VGND VPWR VPWR fd._1580_ sky130_fd_sc_hd__xnor2_1
XFILLER_269_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7392_ fd._2641_ fd._2656_ fd._2657_ VGND VGND VPWR VPWR fd._2658_ sky130_fd_sc_hd__a21o_1
XFILLER_268_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_284_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6343_ fd._1424_ VGND VGND VPWR VPWR fd._1504_ sky130_fd_sc_hd__inv_2
XFILLER_268_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput5 io_in[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6274_ fd._1426_ fd._1423_ fd._1427_ VGND VGND VPWR VPWR fd._1428_ sky130_fd_sc_hd__a21oi_1
XFILLER_133_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_283_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8013_ fd._2076_ fd._3337_ fd._3340_ fd._1330_ VGND VGND VPWR VPWR fd._3341_ sky130_fd_sc_hd__o22ai_1
Xfd._5225_ fd._0273_ fd._0225_ VGND VGND VPWR VPWR fd._0275_ sky130_fd_sc_hd__xnor2_1
XFILLER_188_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5156_ fd._1264_ fd._0073_ fd._0196_ fd._0000_ fd._0198_ VGND VGND VPWR VPWR fd._0199_
+ sky130_fd_sc_hd__a221oi_1
XFILLER_209_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_283_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4107_ fd.a\[0\] fd.b\[0\] VGND VGND VPWR VPWR fd._0362_ sky130_fd_sc_hd__nand2b_1
XFILLER_209_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5087_ fd._3537_ fd._0122_ VGND VGND VPWR VPWR fd._0123_ sky130_fd_sc_hd__xnor2_1
XFILLER_209_1676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_257_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5989_ fd._0946_ fd._1114_ fd._1046_ VGND VGND VPWR VPWR fd._1115_ sky130_fd_sc_hd__mux2_1
XFILLER_203_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7728_ fd._2816_ fd._2819_ VGND VGND VPWR VPWR fd._3028_ sky130_fd_sc_hd__nor2_1
XFILLER_69_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7659_ fd._2751_ fd._2951_ VGND VGND VPWR VPWR fd._2952_ sky130_fd_sc_hd__and2_1
XFILLER_121_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_273_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_262_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_274_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_256_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_282_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_210_ fd.c\[2\] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_1
XFILLER_204_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_254_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_266_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_265_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5010_ fd._3967_ fd._0036_ fd._0037_ VGND VGND VPWR VPWR fd._0038_ sky130_fd_sc_hd__o21a_1
XFILLER_206_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6961_ fd._2179_ fd._2180_ fd._2183_ fd._1976_ VGND VGND VPWR VPWR fd._2184_ sky130_fd_sc_hd__a211o_1
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5912_ fd._0427_ fd._1013_ VGND VGND VPWR VPWR fd._1030_ sky130_fd_sc_hd__nor2_1
XFILLER_187_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6892_ fd._2066_ fd._2104_ fd._2106_ fd._2107_ VGND VGND VPWR VPWR fd._2108_ sky130_fd_sc_hd__o211a_1
XFILLER_35_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5843_ fd._0720_ fd._0898_ fd._0719_ VGND VGND VPWR VPWR fd._0954_ sky130_fd_sc_hd__a21o_1
XFILLER_200_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5774_ fd._0482_ fd._0877_ VGND VGND VPWR VPWR fd._0878_ sky130_fd_sc_hd__nor2_1
XFILLER_192_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7513_ fd._2326_ fd._2790_ VGND VGND VPWR VPWR fd._2791_ sky130_fd_sc_hd__and2_1
XFILLER_115_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4725_ fd._3818_ VGND VGND VPWR VPWR fd._3819_ sky130_fd_sc_hd__clkinv_2
XFILLER_118_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7444_ fd._2517_ fd._2714_ VGND VGND VPWR VPWR fd._2715_ sky130_fd_sc_hd__xnor2_1
XFILLER_135_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4656_ fd._3637_ fd._3748_ fd._3749_ VGND VGND VPWR VPWR fd._3750_ sky130_fd_sc_hd__a21bo_1
XFILLER_29_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_269_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7375_ fd._2433_ fd._2638_ fd._2623_ VGND VGND VPWR VPWR fd._2640_ sky130_fd_sc_hd__mux2_1
Xfd._4587_ fd._3675_ fd._3679_ VGND VGND VPWR VPWR fd._3681_ sky130_fd_sc_hd__nand2_1
XFILLER_170_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_268_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6326_ fd._1483_ fd._1485_ VGND VGND VPWR VPWR fd._1486_ sky130_fd_sc_hd__xnor2_1
XFILLER_111_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_285_1601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_256_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6257_ fd._1409_ VGND VGND VPWR VPWR fd._1410_ sky130_fd_sc_hd__inv_2
XFILLER_168_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5208_ fd._0125_ VGND VGND VPWR VPWR fd._0256_ sky130_fd_sc_hd__inv_2
XFILLER_92_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6188_ fd._0479_ fd._1333_ VGND VGND VPWR VPWR fd._1334_ sky130_fd_sc_hd__nor2_1
XFILLER_240_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_280_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._5139_ fd._0179_ fd._4052_ fd._0060_ VGND VGND VPWR VPWR fd._0180_ sky130_fd_sc_hd__mux2_1
XFILLER_12_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_10 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_268_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_284_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_1612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_9164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_8485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4510_ fd.b\[21\] fd._3603_ VGND VGND VPWR VPWR fd._3604_ sky130_fd_sc_hd__nand2_1
XTAP_7751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_273_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5490_ fd._0292_ fd._0361_ fd._0368_ VGND VGND VPWR VPWR fd._0566_ sky130_fd_sc_hd__a21oi_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_267_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4441_ fd.b\[2\] fd._3534_ VGND VGND VPWR VPWR fd._3535_ sky130_fd_sc_hd__and2_1
XFILLER_39_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_267_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7160_ fd._1656_ fd._2402_ VGND VGND VPWR VPWR fd._2403_ sky130_fd_sc_hd__xnor2_1
XFILLER_43_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_282_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4372_ fd._2441_ fd._3266_ fd._3211_ VGND VGND VPWR VPWR fd._3277_ sky130_fd_sc_hd__mux2_1
XFILLER_226_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6111_ fd._1248_ VGND VGND VPWR VPWR fd._1249_ sky130_fd_sc_hd__inv_2
XFILLER_267_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_253_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7091_ fd._2200_ VGND VGND VPWR VPWR fd._2327_ sky130_fd_sc_hd__clkinv_2
XFILLER_59_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6042_ fd._1172_ VGND VGND VPWR VPWR fd._1173_ sky130_fd_sc_hd__buf_6
XFILLER_130_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_250_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7993_ fd._1102_ fd._3317_ VGND VGND VPWR VPWR fd._3319_ sky130_fd_sc_hd__and2_1
XFILLER_280_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6944_ fd._2142_ fd._2164_ VGND VGND VPWR VPWR fd._2165_ sky130_fd_sc_hd__nor2_1
XFILLER_124_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6875_ fd._2082_ VGND VGND VPWR VPWR fd._2090_ sky130_fd_sc_hd__inv_2
Xinput30 io_in[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_4
XFILLER_50_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5826_ fd._0669_ fd._0676_ fd._0688_ fd._0666_ VGND VGND VPWR VPWR fd._0936_ sky130_fd_sc_hd__a31o_1
XFILLER_85_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5757_ fd._0766_ fd._0859_ fd._0849_ VGND VGND VPWR VPWR fd._0860_ sky130_fd_sc_hd__mux2_1
XFILLER_192_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4708_ fd._3798_ fd._3799_ fd._3800_ fd._3801_ VGND VGND VPWR VPWR fd._3802_ sky130_fd_sc_hd__a31o_1
XFILLER_143_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5688_ fd._0783_ fd._0478_ VGND VGND VPWR VPWR fd._0784_ sky130_fd_sc_hd__xnor2_1
XFILLER_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_269_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4639_ fd._3728_ fd._3731_ fd._3732_ VGND VGND VPWR VPWR fd._3733_ sky130_fd_sc_hd__a21o_1
Xfd._7427_ fd._2604_ fd._2696_ fd._2677_ VGND VGND VPWR VPWR fd._2697_ sky130_fd_sc_hd__mux2_1
XFILLER_285_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_285_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_284_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7358_ fd._2055_ fd._2620_ VGND VGND VPWR VPWR fd._2621_ sky130_fd_sc_hd__xnor2_1
XFILLER_123_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6309_ fd._1459_ fd._1465_ fd._1466_ VGND VGND VPWR VPWR fd._1467_ sky130_fd_sc_hd__a21oi_1
Xfd._7289_ fd._2376_ fd._2379_ VGND VGND VPWR VPWR fd._2545_ sky130_fd_sc_hd__or2_1
XFILLER_42_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_285_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1531 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_249_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1580 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_264_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_264_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._4990_ fd._3972_ fd._0008_ fd._0014_ fd._0015_ VGND VGND VPWR VPWR fd._0016_ sky130_fd_sc_hd__a31oi_2
XFILLER_121_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6660_ fd._1851_ VGND VGND VPWR VPWR fd._1853_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_8_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5611_ fd._0697_ fd._0666_ fd._0695_ VGND VGND VPWR VPWR fd._0699_ sky130_fd_sc_hd__o21a_1
XFILLER_67_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6591_ fd._0928_ fd._1735_ VGND VGND VPWR VPWR fd._1777_ sky130_fd_sc_hd__nand2_1
XFILLER_171_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_275_1699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5542_ fd._0450_ fd._0622_ VGND VGND VPWR VPWR fd._0623_ sky130_fd_sc_hd__xnor2_1
XFILLER_125_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._8261_ net70 net14 VGND VGND VPWR VPWR fd.b\[21\] sky130_fd_sc_hd__dfxtp_2
XTAP_7592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5473_ fd._0541_ fd._0546_ VGND VGND VPWR VPWR fd._0547_ sky130_fd_sc_hd__nor2_1
XFILLER_6_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7212_ fd._2427_ fd._2433_ VGND VGND VPWR VPWR fd._2460_ sky130_fd_sc_hd__or2_1
XFILLER_266_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4424_ fd._3515_ fd._3517_ VGND VGND VPWR VPWR fd._3518_ sky130_fd_sc_hd__xor2_1
XTAP_6891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._8192_ net71 fd.mc\[16\] VGND VGND VPWR VPWR fd.c\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_267_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7143_ fd._1751_ fd._2366_ VGND VGND VPWR VPWR fd._2384_ sky130_fd_sc_hd__nor2_1
XFILLER_282_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4355_ fd._1132_ fd._3079_ VGND VGND VPWR VPWR fd._3090_ sky130_fd_sc_hd__or2_1
XFILLER_26_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7074_ fd._1242_ fd._2307_ VGND VGND VPWR VPWR fd._2308_ sky130_fd_sc_hd__or2_1
Xfd._4286_ fd._1572_ fd._1616_ VGND VGND VPWR VPWR fd._2331_ sky130_fd_sc_hd__nand2_1
XFILLER_235_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6025_ fd._1275_ fd._1152_ VGND VGND VPWR VPWR fd._1155_ sky130_fd_sc_hd__and2_1
XFILLER_34_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7976_ fd._3149_ fd._3300_ VGND VGND VPWR VPWR fd._3301_ sky130_fd_sc_hd__xnor2_1
Xfd._6927_ fd._1949_ fd._1984_ VGND VGND VPWR VPWR fd._2147_ sky130_fd_sc_hd__and2b_1
XFILLER_163_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6858_ fd._2068_ fd._2070_ VGND VGND VPWR VPWR fd._2071_ sky130_fd_sc_hd__xnor2_1
XFILLER_116_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_254_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5809_ fd._0916_ fd._0914_ VGND VGND VPWR VPWR fd._0917_ sky130_fd_sc_hd__and2_1
XFILLER_150_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6789_ fd._1173_ fd._1930_ VGND VGND VPWR VPWR fd._1995_ sky130_fd_sc_hd__or2_1
XFILLER_143_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_1548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_285_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_214_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_279_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_279_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_208 VGND VGND VPWR VPWR user_project_wrapper_208/HI la_data_out[86]
+ sky130_fd_sc_hd__conb_1
XFILLER_153_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_219 VGND VGND VPWR VPWR user_project_wrapper_219/HI la_data_out[97]
+ sky130_fd_sc_hd__conb_1
XFILLER_119_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_1604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4140_ fd._0681_ fd._0714_ VGND VGND VPWR VPWR fd._0725_ sky130_fd_sc_hd__nand2_1
XTAP_4796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_251_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_262_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._7830_ fd._2135_ fd._3139_ VGND VGND VPWR VPWR fd._3140_ sky130_fd_sc_hd__nor2_1
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4973_ fd._1297_ fd._4067_ VGND VGND VPWR VPWR fd._4069_ sky130_fd_sc_hd__nand2_1
Xfd._7761_ fd._3063_ fd._3062_ VGND VGND VPWR VPWR fd._3064_ sky130_fd_sc_hd__nor2_1
XFILLER_258_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6712_ fd._1632_ fd._1828_ VGND VGND VPWR VPWR fd._1910_ sky130_fd_sc_hd__nor2_1
XFILLER_51_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7692_ fd._2977_ fd._2984_ fd._2986_ fd._2987_ VGND VGND VPWR VPWR fd._2988_ sky130_fd_sc_hd__a211o_1
XFILLER_12_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6643_ fd._1165_ fd._1823_ VGND VGND VPWR VPWR fd._1834_ sky130_fd_sc_hd__nor2_1
XFILLER_132_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6574_ fd._1757_ fd._1589_ VGND VGND VPWR VPWR fd._1758_ sky130_fd_sc_hd__or2_1
XFILLER_119_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5525_ fd._0392_ fd._0603_ fd._0453_ VGND VGND VPWR VPWR fd._0605_ sky130_fd_sc_hd__mux2_1
XFILLER_119_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_269_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8244_ net72 net27 VGND VGND VPWR VPWR fd.b\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_228_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5456_ fd._0311_ fd._0528_ VGND VGND VPWR VPWR fd._0529_ sky130_fd_sc_hd__xnor2_1
XFILLER_230_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4407_ fd._3499_ fd._3500_ VGND VGND VPWR VPWR fd._3501_ sky130_fd_sc_hd__xnor2_1
XFILLER_254_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8175_ fd.b\[31\] fd.a\[31\] VGND VGND VPWR VPWR fd.sc sky130_fd_sc_hd__xor2_1
XFILLER_66_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5387_ fd._0452_ VGND VGND VPWR VPWR fd._0453_ sky130_fd_sc_hd__buf_6
XFILLER_82_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7126_ fd._2173_ fd._2365_ fd._2322_ VGND VGND VPWR VPWR fd._2366_ sky130_fd_sc_hd__mux2_1
Xfd._4338_ fd._1055_ fd._2848_ VGND VGND VPWR VPWR fd._2903_ sky130_fd_sc_hd__xnor2_1
XFILLER_270_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_247_1543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7057_ fd._2284_ fd._2288_ fd._2289_ VGND VGND VPWR VPWR fd._2290_ sky130_fd_sc_hd__o21bai_1
XFILLER_78_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4269_ fd._1704_ fd._2078_ fd._2122_ fd._2133_ VGND VGND VPWR VPWR fd._2144_ sky130_fd_sc_hd__o31a_1
XFILLER_35_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6008_ fd._1134_ fd._1135_ VGND VGND VPWR VPWR fd._1136_ sky130_fd_sc_hd__nor2_1
XFILLER_223_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7959_ fd._3169_ fd._3171_ fd._3172_ VGND VGND VPWR VPWR fd._3282_ sky130_fd_sc_hd__a21o_1
XFILLER_175_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_277_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_1663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_268_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_283_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5310_ fd._0365_ fd._0367_ VGND VGND VPWR VPWR fd._0368_ sky130_fd_sc_hd__nor2_1
XFILLER_7_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6290_ fd._1274_ fd._1273_ VGND VGND VPWR VPWR fd._1446_ sky130_fd_sc_hd__or2b_1
XTAP_5250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_283_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5241_ fd._3833_ fd._0291_ VGND VGND VPWR VPWR fd._0292_ sky130_fd_sc_hd__or2_1
XTAP_5283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_266_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5172_ fd._0026_ fd._0214_ VGND VGND VPWR VPWR fd._0216_ sky130_fd_sc_hd__and2_1
XFILLER_221_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4123_ fd.a\[9\] VGND VGND VPWR VPWR fd._0538_ sky130_fd_sc_hd__inv_2
XFILLER_252_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_251_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7813_ fd._3119_ fd._3120_ VGND VGND VPWR VPWR fd._3121_ sky130_fd_sc_hd__nand2_1
XFILLER_121_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7744_ fd._3029_ fd._2839_ VGND VGND VPWR VPWR fd._3045_ sky130_fd_sc_hd__xor2_1
XFILLER_121_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4956_ fd._3917_ fd._4050_ VGND VGND VPWR VPWR fd._4051_ sky130_fd_sc_hd__or2_1
XFILLER_195_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4887_ fd._3469_ fd._3975_ fd._3979_ fd._3980_ VGND VGND VPWR VPWR fd._3981_ sky130_fd_sc_hd__o22a_1
XFILLER_195_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7675_ fd._2966_ fd._2876_ fd._2967_ fd._2968_ VGND VGND VPWR VPWR fd._2970_ sky130_fd_sc_hd__o31a_1
XFILLER_133_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6626_ fd._0786_ VGND VGND VPWR VPWR fd._1816_ sky130_fd_sc_hd__buf_6
XFILLER_132_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6557_ fd._1566_ VGND VGND VPWR VPWR fd._1740_ sky130_fd_sc_hd__inv_2
XFILLER_59_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5508_ fd._0375_ fd._0379_ fd._0385_ VGND VGND VPWR VPWR fd._0586_ sky130_fd_sc_hd__a21oi_1
XFILLER_189_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6488_ fd._1448_ fd._1663_ fd._1615_ VGND VGND VPWR VPWR fd._1664_ sky130_fd_sc_hd__mux2_1
XFILLER_101_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_1586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8227_ net70 net11 VGND VGND VPWR VPWR fd.a\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_255_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5439_ fd._0508_ fd._0509_ VGND VGND VPWR VPWR fd._0510_ sky130_fd_sc_hd__xnor2_1
XFILLER_67_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8158_ fd._3466_ fd._3472_ VGND VGND VPWR VPWR fd._3473_ sky130_fd_sc_hd__nor2_1
XFILLER_83_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7109_ fd._2339_ fd._2345_ fd._2346_ VGND VGND VPWR VPWR fd._2347_ sky130_fd_sc_hd__a21oi_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8089_ fd._1232_ fd._1423_ fd._3411_ VGND VGND VPWR VPWR fd._3413_ sky130_fd_sc_hd__mux2_1
XFILLER_224_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_282_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_265_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_283_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_281_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_259_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._4810_ fd._0857_ fd._3903_ VGND VGND VPWR VPWR fd._3904_ sky130_fd_sc_hd__and2_1
Xfd._5790_ fd._0726_ fd._0894_ VGND VGND VPWR VPWR fd._0896_ sky130_fd_sc_hd__nor2_1
XFILLER_128_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_1545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4741_ fd._3716_ fd._3720_ VGND VGND VPWR VPWR fd._3835_ sky130_fd_sc_hd__and2_1
XFILLER_202_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4672_ fd._3603_ fd._3765_ fd._3626_ VGND VGND VPWR VPWR fd._3766_ sky130_fd_sc_hd__mux2_1
Xfd._7460_ fd._2730_ fd._2732_ VGND VGND VPWR VPWR fd._2733_ sky130_fd_sc_hd__xnor2_1
XFILLER_272_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6411_ fd._1578_ fd._1398_ VGND VGND VPWR VPWR fd._1579_ sky130_fd_sc_hd__and2b_1
Xfd._7391_ fd._2481_ fd._2635_ VGND VGND VPWR VPWR fd._2657_ sky130_fd_sc_hd__xnor2_1
XFILLER_123_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6342_ fd._1434_ fd._1500_ fd._1502_ VGND VGND VPWR VPWR fd._1503_ sky130_fd_sc_hd__a21o_1
XFILLER_155_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6273_ fd._1301_ fd._1340_ fd._1348_ VGND VGND VPWR VPWR fd._1427_ sky130_fd_sc_hd__and3_1
Xinput6 io_in[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5224_ fd._0272_ fd._0218_ fd._0215_ VGND VGND VPWR VPWR fd._0273_ sky130_fd_sc_hd__a21oi_1
Xfd._8012_ fd._3102_ fd._3339_ fd._3240_ VGND VGND VPWR VPWR fd._3340_ sky130_fd_sc_hd__mux2_1
XFILLER_237_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5155_ fd._0190_ fd._0194_ VGND VGND VPWR VPWR fd._0198_ sky130_fd_sc_hd__nor2_1
XFILLER_206_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4106_ fd._0329_ fd._0340_ VGND VGND VPWR VPWR fd._0351_ sky130_fd_sc_hd__nor2_1
XFILLER_33_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5086_ fd._3695_ fd._3961_ VGND VGND VPWR VPWR fd._0122_ sky130_fd_sc_hd__nor2_1
XFILLER_209_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5988_ fd._0942_ fd._1113_ VGND VGND VPWR VPWR fd._1114_ sky130_fd_sc_hd__xnor2_1
XFILLER_134_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7727_ fd._2843_ VGND VGND VPWR VPWR fd._3027_ sky130_fd_sc_hd__inv_2
Xfd._4939_ fd._0868_ fd._4032_ VGND VGND VPWR VPWR fd._4033_ sky130_fd_sc_hd__nand2_1
XFILLER_118_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7658_ fd._2945_ fd._2950_ fd._2874_ VGND VGND VPWR VPWR fd._2951_ sky130_fd_sc_hd__mux2_1
XFILLER_82_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6609_ fd._0541_ VGND VGND VPWR VPWR fd._1797_ sky130_fd_sc_hd__buf_6
XFILLER_173_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_1659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7589_ fd._2874_ VGND VGND VPWR VPWR fd._2875_ sky130_fd_sc_hd__buf_8
XFILLER_113_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_256_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_255_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_271_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_282_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1635 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_9313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_267_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_265_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_261_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_1506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._6960_ fd._2033_ fd._2048_ fd._2113_ fd._2182_ VGND VGND VPWR VPWR fd._2183_ sky130_fd_sc_hd__o31a_1
XFILLER_124_1517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._5911_ fd._1015_ fd._1019_ fd._1025_ fd._1028_ VGND VGND VPWR VPWR fd._1029_ sky130_fd_sc_hd__o211ai_2
XFILLER_147_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6891_ fd._0207_ fd._2061_ VGND VGND VPWR VPWR fd._2107_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5842_ fd._0903_ fd._0952_ fd._3917_ VGND VGND VPWR VPWR fd._0953_ sky130_fd_sc_hd__a21o_1
XFILLER_278_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5773_ fd._0755_ fd._0875_ fd._0849_ fd._0876_ VGND VGND VPWR VPWR fd._0877_ sky130_fd_sc_hd__a31oi_4
XFILLER_196_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7512_ fd._2787_ fd._2789_ fd._2677_ VGND VGND VPWR VPWR fd._2790_ sky130_fd_sc_hd__mux2_1
XFILLER_48_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4724_ fd._3733_ fd._3737_ VGND VGND VPWR VPWR fd._3818_ sky130_fd_sc_hd__xnor2_1
XFILLER_142_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_1640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7443_ fd._2523_ fd._2565_ VGND VGND VPWR VPWR fd._2714_ sky130_fd_sc_hd__and2_1
Xfd._4655_ fd._3580_ fd._3632_ VGND VGND VPWR VPWR fd._3749_ sky130_fd_sc_hd__nand2_1
XFILLER_233_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_272_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_269_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4586_ fd._3675_ fd._3679_ VGND VGND VPWR VPWR fd._3680_ sky130_fd_sc_hd__or2_1
XFILLER_233_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7374_ fd._2462_ fd._2637_ VGND VGND VPWR VPWR fd._2638_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6325_ fd._1241_ fd._1282_ VGND VGND VPWR VPWR fd._1485_ sky130_fd_sc_hd__and2_1
XFILLER_238_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_284_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6256_ fd._1183_ fd._1408_ fd._1349_ VGND VGND VPWR VPWR fd._1409_ sky130_fd_sc_hd__mux2_1
XFILLER_42_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_271_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_253_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5207_ fd._0242_ fd._0244_ fd._0254_ fd._0246_ VGND VGND VPWR VPWR fd._0255_ sky130_fd_sc_hd__a22o_1
XFILLER_227_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6187_ fd._1332_ VGND VGND VPWR VPWR fd._1333_ sky130_fd_sc_hd__inv_2
XFILLER_52_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5138_ fd._4047_ fd._0178_ VGND VGND VPWR VPWR fd._0179_ sky130_fd_sc_hd__xnor2_1
XFILLER_52_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5069_ fd._0102_ fd._3998_ fd._0059_ VGND VGND VPWR VPWR fd._0103_ sky130_fd_sc_hd__mux2_1
XFILLER_178_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_11 fd._1644_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_1641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_268_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_255_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_251_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_251_1358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_8464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4440_ fd._3523_ fd._3533_ fd._3200_ VGND VGND VPWR VPWR fd._3534_ sky130_fd_sc_hd__mux2_1
XTAP_7796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_267_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_1578 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4371_ fd._3255_ VGND VGND VPWR VPWR fd._3266_ sky130_fd_sc_hd__clkinv_2
XFILLER_117_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_266_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_282_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6110_ fd._1246_ fd._1247_ VGND VGND VPWR VPWR fd._1248_ sky130_fd_sc_hd__and2_1
XFILLER_47_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7090_ fd._0343_ VGND VGND VPWR VPWR fd._2326_ sky130_fd_sc_hd__buf_6
XFILLER_267_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_281_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6041_ fd._0662_ VGND VGND VPWR VPWR fd._1172_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_185_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_267_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_261_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_280_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7992_ fd._1797_ fd._3313_ fd._3317_ fd._1102_ VGND VGND VPWR VPWR fd._3318_ sky130_fd_sc_hd__o22ai_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6943_ fd._2159_ fd._2163_ fd._2115_ VGND VGND VPWR VPWR fd._2164_ sky130_fd_sc_hd__mux2_1
XFILLER_124_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput20 io_in[27] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_1
XFILLER_204_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6874_ fd._1118_ fd._2087_ VGND VGND VPWR VPWR fd._2088_ sky130_fd_sc_hd__nor2_1
Xinput31 io_in[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_4
XFILLER_239_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5825_ fd._0919_ fd._0925_ fd._0927_ fd._0930_ fd._0933_ VGND VGND VPWR VPWR fd._0935_
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_239_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5756_ fd._0851_ fd._0852_ VGND VGND VPWR VPWR fd._0859_ sky130_fd_sc_hd__xnor2_1
XFILLER_157_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_1601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_277_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4707_ fd._3632_ fd._3788_ VGND VGND VPWR VPWR fd._3801_ sky130_fd_sc_hd__and2_1
XFILLER_153_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5687_ fd._0469_ fd._0782_ fd._0480_ VGND VGND VPWR VPWR fd._0783_ sky130_fd_sc_hd__o21a_1
XFILLER_258_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7426_ fd._2601_ fd._2695_ VGND VGND VPWR VPWR fd._2696_ sky130_fd_sc_hd__xnor2_1
Xfd._4638_ fd.b\[13\] fd._3730_ VGND VGND VPWR VPWR fd._3732_ sky130_fd_sc_hd__and2_1
XFILLER_229_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_285_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7357_ fd._2618_ fd._2619_ fd._2506_ VGND VGND VPWR VPWR fd._2620_ sky130_fd_sc_hd__mux2_1
Xfd._4569_ fd._3662_ VGND VGND VPWR VPWR fd._3663_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_245_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_268_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6308_ fd._0846_ fd._1464_ VGND VGND VPWR VPWR fd._1466_ sky130_fd_sc_hd__nor2_1
XFILLER_84_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7288_ fd._2142_ fd._2543_ VGND VGND VPWR VPWR fd._2544_ sky130_fd_sc_hd__xnor2_1
XFILLER_272_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6239_ fd._1015_ fd._1389_ VGND VGND VPWR VPWR fd._1390_ sky130_fd_sc_hd__nand2_1
XFILLER_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_279_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_279_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_257_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_1507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_249_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_249_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_251_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_272_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5610_ fd._0696_ fd._0697_ VGND VGND VPWR VPWR fd._0698_ sky130_fd_sc_hd__nor2_1
XFILLER_271_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_8250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._6590_ fd._1756_ fd._1762_ fd._1773_ fd._1774_ fd._1775_ VGND VGND VPWR VPWR fd._1776_
+ sky130_fd_sc_hd__o311a_1
XFILLER_67_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_259_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5541_ fd._0435_ fd._0621_ fd._0613_ VGND VGND VPWR VPWR fd._0622_ sky130_fd_sc_hd__mux2_1
XFILLER_3_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8260_ net70 net13 VGND VGND VPWR VPWR fd.b\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_7582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5472_ fd._0542_ fd._0545_ fd._0452_ VGND VGND VPWR VPWR fd._0546_ sky130_fd_sc_hd__mux2_1
XFILLER_39_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7211_ fd._1494_ fd._2439_ fd._2453_ fd._2458_ VGND VGND VPWR VPWR fd._2459_ sky130_fd_sc_hd__a31o_1
XFILLER_45_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4423_ fd._1891_ fd._3516_ VGND VGND VPWR VPWR fd._3517_ sky130_fd_sc_hd__nand2_1
XTAP_6892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8191_ net73 fd.mc\[15\] VGND VGND VPWR VPWR fd.c\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_227_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4354_ fd._0175_ fd._1077_ fd._1121_ VGND VGND VPWR VPWR fd._3079_ sky130_fd_sc_hd__and3_1
Xfd._7142_ fd._1958_ fd._2373_ fd._2380_ fd._2382_ VGND VGND VPWR VPWR fd._2383_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_43_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_254_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4285_ fd._2144_ fd._2221_ fd._2298_ fd._2309_ VGND VGND VPWR VPWR fd._2320_ sky130_fd_sc_hd__o31a_1
Xfd._7073_ fd._2041_ fd._2238_ fd._2306_ VGND VGND VPWR VPWR fd._2307_ sky130_fd_sc_hd__o21a_1
XFILLER_81_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6024_ fd._1275_ fd._1152_ VGND VGND VPWR VPWR fd._1153_ sky130_fd_sc_hd__or2_1
XFILLER_78_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_222_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_280_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7975_ fd._3152_ fd._3177_ VGND VGND VPWR VPWR fd._3300_ sky130_fd_sc_hd__nor2_1
XFILLER_187_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6926_ fd._2143_ fd._2145_ fd._1983_ VGND VGND VPWR VPWR fd._2146_ sky130_fd_sc_hd__a21bo_1
XFILLER_50_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6857_ fd._2069_ fd._1895_ VGND VGND VPWR VPWR fd._2070_ sky130_fd_sc_hd__nor2_1
XFILLER_50_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5808_ fd._0089_ VGND VGND VPWR VPWR fd._0916_ sky130_fd_sc_hd__buf_6
XFILLER_11_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6788_ fd._0928_ fd._1989_ VGND VGND VPWR VPWR fd._1994_ sky130_fd_sc_hd__nor2_1
XFILLER_89_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5739_ fd._0775_ fd._0795_ fd._0781_ VGND VGND VPWR VPWR fd._0840_ sky130_fd_sc_hd__a21o_1
XFILLER_172_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_277_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_1551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7409_ fd._2676_ VGND VGND VPWR VPWR fd._2677_ sky130_fd_sc_hd__buf_8
XTAP_4208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_272_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_279_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_279_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_project_wrapper_209 VGND VGND VPWR VPWR user_project_wrapper_209/HI la_data_out[87]
+ sky130_fd_sc_hd__conb_1
XFILLER_111_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_1586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_264_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_249_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_1543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7760_ fd._3019_ fd._3020_ VGND VGND VPWR VPWR fd._3063_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4972_ fd._1297_ fd._4067_ VGND VGND VPWR VPWR fd._4068_ sky130_fd_sc_hd__or2_1
XFILLER_219_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6711_ fd._1632_ fd._1828_ VGND VGND VPWR VPWR fd._1909_ sky130_fd_sc_hd__and2_1
XFILLER_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7691_ fd._1656_ fd._2983_ VGND VGND VPWR VPWR fd._2987_ sky130_fd_sc_hd__nor2_1
XFILLER_12_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6642_ fd._1815_ fd._1832_ VGND VGND VPWR VPWR fd._1833_ sky130_fd_sc_hd__nand2_1
XFILLER_12_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1448 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_259_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._6573_ fd._1397_ fd._1588_ VGND VGND VPWR VPWR fd._1757_ sky130_fd_sc_hd__nor2_1
XFILLER_4_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5524_ fd._0397_ fd._0602_ VGND VGND VPWR VPWR fd._0603_ sky130_fd_sc_hd__nand2_1
XFILLER_141_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_1402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8243_ net74 net26 VGND VGND VPWR VPWR fd.b\[3\] sky130_fd_sc_hd__dfxtp_2
XFILLER_267_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5455_ fd._0317_ fd._0328_ VGND VGND VPWR VPWR fd._0528_ sky130_fd_sc_hd__or2_1
XFILLER_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4406_ fd._1704_ fd._2067_ VGND VGND VPWR VPWR fd._3500_ sky130_fd_sc_hd__or2_1
XFILLER_132_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_282_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8174_ fd._3483_ fd._3487_ VGND VGND VPWR VPWR fd.ec\[7\] sky130_fd_sc_hd__xnor2_1
XFILLER_254_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5386_ fd._0425_ VGND VGND VPWR VPWR fd._0452_ sky130_fd_sc_hd__buf_6
XFILLER_269_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7125_ fd._2361_ fd._2363_ VGND VGND VPWR VPWR fd._2365_ sky130_fd_sc_hd__xnor2_1
XFILLER_81_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4337_ fd.b\[20\] fd._2881_ VGND VGND VPWR VPWR fd._2892_ sky130_fd_sc_hd__or2_1
XFILLER_254_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7056_ fd._1275_ fd._2260_ VGND VGND VPWR VPWR fd._2289_ sky130_fd_sc_hd__nor2_1
XFILLER_39_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4268_ fd._0428_ fd._2111_ VGND VGND VPWR VPWR fd._2133_ sky130_fd_sc_hd__or2_1
XFILLER_251_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6007_ fd._0953_ fd._0959_ fd._0897_ VGND VGND VPWR VPWR fd._1135_ sky130_fd_sc_hd__a21oi_1
XFILLER_180_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4199_ fd._1363_ fd._1000_ VGND VGND VPWR VPWR fd._1374_ sky130_fd_sc_hd__xnor2_1
XFILLER_195_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7958_ fd._2751_ fd._3267_ fd._3270_ fd._3280_ VGND VGND VPWR VPWR fd._3281_ sky130_fd_sc_hd__o211a_1
XFILLER_30_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_276_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6909_ fd._1994_ fd._1991_ VGND VGND VPWR VPWR fd._2127_ sky130_fd_sc_hd__and2b_1
XFILLER_190_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7889_ fd._3096_ fd._3204_ VGND VGND VPWR VPWR fd._3205_ sky130_fd_sc_hd__and2_1
XFILLER_135_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_1330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5240_ fd._0161_ fd._0290_ fd._0269_ VGND VGND VPWR VPWR fd._0291_ sky130_fd_sc_hd__mux2_1
XTAP_5273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5171_ fd._0026_ fd._0214_ VGND VGND VPWR VPWR fd._0215_ sky130_fd_sc_hd__nor2_1
XTAP_4583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4122_ fd.b\[9\] fd.a\[9\] VGND VGND VPWR VPWR fd._0527_ sky130_fd_sc_hd__nand2b_1
XTAP_3882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_233_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_260_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_1463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7812_ fd._3104_ fd._3099_ VGND VGND VPWR VPWR fd._3120_ sky130_fd_sc_hd__and2b_1
XFILLER_242_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_277_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7743_ fd._2835_ VGND VGND VPWR VPWR fd._3044_ sky130_fd_sc_hd__clkinv_2
Xfd._4955_ fd._3838_ fd._4048_ fd._3960_ VGND VGND VPWR VPWR fd._4050_ sky130_fd_sc_hd__mux2_1
XFILLER_172_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7674_ fd._2734_ fd._2876_ VGND VGND VPWR VPWR fd._2968_ sky130_fd_sc_hd__nand2_1
Xfd._4886_ fd._2155_ VGND VGND VPWR VPWR fd._3980_ sky130_fd_sc_hd__buf_6
XFILLER_172_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6625_ fd._1639_ fd._1812_ fd._1813_ VGND VGND VPWR VPWR fd._1815_ sky130_fd_sc_hd__mux2_2
XFILLER_173_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6556_ fd._1574_ fd._1593_ fd._1573_ VGND VGND VPWR VPWR fd._1739_ sky130_fd_sc_hd__a21oi_1
XFILLER_119_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5507_ fd._0579_ fd._0967_ fd._0584_ VGND VGND VPWR VPWR fd._0585_ sky130_fd_sc_hd__mux2_1
XFILLER_268_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6487_ fd._0716_ fd._1468_ VGND VGND VPWR VPWR fd._1663_ sky130_fd_sc_hd__xnor2_1
XFILLER_140_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8226_ net70 net10 VGND VGND VPWR VPWR fd.a\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_269_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5438_ fd._0317_ fd._0326_ VGND VGND VPWR VPWR fd._0509_ sky130_fd_sc_hd__or2b_1
XFILLER_210_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_255_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_270_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8157_ fd._3470_ fd._3471_ VGND VGND VPWR VPWR fd._3472_ sky130_fd_sc_hd__nor2_1
XFILLER_82_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5369_ fd._0432_ fd._0257_ VGND VGND VPWR VPWR fd._0433_ sky130_fd_sc_hd__nor2_1
XFILLER_215_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7108_ fd._1600_ fd._2338_ VGND VGND VPWR VPWR fd._2346_ sky130_fd_sc_hd__and2_1
XFILLER_36_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8088_ fd._3412_ VGND VGND VPWR VPWR fd.mc\[11\] sky130_fd_sc_hd__clkbuf_1
XFILLER_184_1631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7039_ fd._2223_ fd._2227_ fd._2269_ fd._2267_ VGND VGND VPWR VPWR fd._2270_ sky130_fd_sc_hd__a31o_1
XFILLER_24_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_1528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_260_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_8838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_246_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_259_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4740_ fd._3651_ fd._3715_ VGND VGND VPWR VPWR fd._3834_ sky130_fd_sc_hd__or2_1
XFILLER_155_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_259_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4671_ fd._3606_ fd._3764_ VGND VGND VPWR VPWR fd._3765_ sky130_fd_sc_hd__xnor2_1
XFILLER_29_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6410_ fd._1397_ fd._1576_ VGND VGND VPWR VPWR fd._1578_ sky130_fd_sc_hd__nor2_1
XFILLER_116_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_268_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7390_ fd._2645_ fd._2654_ fd._2655_ VGND VGND VPWR VPWR fd._2656_ sky130_fd_sc_hd__a21bo_1
XFILLER_237_1598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6341_ fd._1430_ fd._1501_ VGND VGND VPWR VPWR fd._1502_ sky130_fd_sc_hd__nand2_1
XFILLER_268_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6272_ fd._1302_ fd._1298_ VGND VGND VPWR VPWR fd._1426_ sky130_fd_sc_hd__xnor2_1
XTAP_5070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput7 io_in[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_237_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._8011_ fd._3119_ fd._3338_ VGND VGND VPWR VPWR fd._3339_ sky130_fd_sc_hd__xnor2_1
XFILLER_65_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_266_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5223_ fd._0070_ fd._0211_ VGND VGND VPWR VPWR fd._0272_ sky130_fd_sc_hd__and2_1
XFILLER_265_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5154_ fd._0190_ fd._0195_ VGND VGND VPWR VPWR fd._0196_ sky130_fd_sc_hd__xnor2_1
XFILLER_209_1601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_252_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4105_ fd.a\[2\] fd.b\[2\] VGND VGND VPWR VPWR fd._0340_ sky130_fd_sc_hd__and2b_1
XFILLER_209_1634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5085_ fd._3689_ fd._3961_ VGND VGND VPWR VPWR fd._0121_ sky130_fd_sc_hd__nand2_1
XFILLER_221_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_257_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5987_ fd._0950_ fd._0947_ VGND VGND VPWR VPWR fd._1113_ sky130_fd_sc_hd__nand2_1
XFILLER_195_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_277_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7726_ fd._2861_ fd._3025_ fd._2877_ VGND VGND VPWR VPWR fd._3026_ sky130_fd_sc_hd__mux2_1
XFILLER_134_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4938_ fd._4029_ fd._4031_ fd._3960_ VGND VGND VPWR VPWR fd._4032_ sky130_fd_sc_hd__mux2_1
XFILLER_133_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7657_ fd._2946_ fd._2949_ VGND VGND VPWR VPWR fd._2950_ sky130_fd_sc_hd__xnor2_1
XFILLER_133_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4869_ fd._3962_ VGND VGND VPWR VPWR fd._3963_ sky130_fd_sc_hd__inv_2
XFILLER_195_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6608_ fd._1788_ fd._1794_ fd._1795_ VGND VGND VPWR VPWR fd._1796_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7588_ fd._2851_ fd._2866_ fd._2868_ fd._2873_ VGND VGND VPWR VPWR fd._2874_ sky130_fd_sc_hd__a211o_4
XFILLER_59_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_275_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._6539_ fd._1719_ VGND VGND VPWR VPWR fd._1720_ sky130_fd_sc_hd__buf_6
XFILLER_19_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8209_ net74 net12 VGND VGND VPWR VPWR fd.a\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_27_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_282_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_1590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_279_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_265_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_281_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5910_ fd._0638_ fd._1026_ fd._1027_ fd._0632_ VGND VGND VPWR VPWR fd._1028_ sky130_fd_sc_hd__a211o_1
XFILLER_41_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6890_ fd._2054_ fd._2105_ VGND VGND VPWR VPWR fd._2106_ sky130_fd_sc_hd__nor2_1
XFILLER_30_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5841_ fd._0942_ fd._0947_ fd._0949_ fd._0951_ VGND VGND VPWR VPWR fd._0952_ sky130_fd_sc_hd__a211o_1
XFILLER_196_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5772_ fd._0753_ fd._0849_ VGND VGND VPWR VPWR fd._0876_ sky130_fd_sc_hd__nor2_1
XFILLER_196_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7511_ fd._2788_ fd._2574_ VGND VGND VPWR VPWR fd._2789_ sky130_fd_sc_hd__xor2_1
Xfd._4723_ fd._2584_ fd._3816_ VGND VGND VPWR VPWR fd._3817_ sky130_fd_sc_hd__nand2_1
XFILLER_170_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_272_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7442_ fd._2712_ VGND VGND VPWR VPWR fd._2713_ sky130_fd_sc_hd__inv_2
Xfd._4654_ fd._3645_ fd._3745_ fd._3747_ VGND VGND VPWR VPWR fd._3748_ sky130_fd_sc_hd__a21o_1
XFILLER_130_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._7373_ fd._2454_ fd._2459_ VGND VGND VPWR VPWR fd._2637_ sky130_fd_sc_hd__nand2_1
XFILLER_116_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4585_ fd._3530_ fd._3678_ fd._3624_ VGND VGND VPWR VPWR fd._3679_ sky130_fd_sc_hd__mux2_1
XFILLER_110_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_284_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6324_ fd._1278_ fd._1281_ VGND VGND VPWR VPWR fd._1483_ sky130_fd_sc_hd__or2_1
XFILLER_81_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_250_1573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_285_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6255_ fd._1185_ fd._1406_ VGND VGND VPWR VPWR fd._1408_ sky130_fd_sc_hd__xnor2_1
XFILLER_49_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_266_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5206_ fd._4011_ fd._0129_ VGND VGND VPWR VPWR fd._0254_ sky130_fd_sc_hd__nand2_1
XFILLER_20_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6186_ fd._1068_ fd._1331_ fd._1232_ VGND VGND VPWR VPWR fd._1332_ sky130_fd_sc_hd__mux2_1
XFILLER_65_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5137_ fd._4053_ fd._4051_ VGND VGND VPWR VPWR fd._0178_ sky130_fd_sc_hd__and2b_1
XFILLER_94_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_283_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5068_ fd._0092_ fd._0101_ VGND VGND VPWR VPWR fd._0102_ sky130_fd_sc_hd__nand2_1
XFILLER_181_1656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_12 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7709_ fd._0382_ fd._3005_ VGND VGND VPWR VPWR fd._3007_ sky130_fd_sc_hd__nand2_1
XFILLER_12_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_262_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_249_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1663 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_256_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_1669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_266_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4370_ fd._3244_ fd._2485_ VGND VGND VPWR VPWR fd._3255_ sky130_fd_sc_hd__xor2_1
XFILLER_94_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6040_ fd._1170_ VGND VGND VPWR VPWR fd._1171_ sky130_fd_sc_hd__clkinv_2
XFILLER_130_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_250_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7991_ fd._3183_ fd._3316_ fd._3239_ VGND VGND VPWR VPWR fd._3317_ sky130_fd_sc_hd__mux2_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._6942_ fd._2160_ fd._2162_ VGND VGND VPWR VPWR fd._2163_ sky130_fd_sc_hd__xor2_1
XFILLER_230_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput10 io_in[18] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_200_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6873_ fd._1877_ fd._2086_ fd._1917_ VGND VGND VPWR VPWR fd._2087_ sky130_fd_sc_hd__mux2_1
XFILLER_147_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput21 io_in[28] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_1
XFILLER_163_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput32 io_in[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_2
XFILLER_156_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5824_ fd._0932_ VGND VGND VPWR VPWR fd._0933_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_50_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5755_ fd._0843_ fd._0844_ fd._0850_ fd._0856_ VGND VGND VPWR VPWR fd._0858_ sky130_fd_sc_hd__o22a_2
XFILLER_171_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1700 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4706_ fd._3787_ VGND VGND VPWR VPWR fd._3800_ sky130_fd_sc_hd__clkinv_8
XFILLER_170_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5686_ fd._0772_ fd._0608_ fd._0476_ VGND VGND VPWR VPWR fd._0782_ sky130_fd_sc_hd__o21bai_1
XFILLER_83_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_276_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_269_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7425_ fd._2607_ fd._2693_ VGND VGND VPWR VPWR fd._2695_ sky130_fd_sc_hd__nand2_1
XFILLER_48_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4637_ fd.b\[13\] fd._3730_ VGND VGND VPWR VPWR fd._3731_ sky130_fd_sc_hd__or2_1
XFILLER_252_1668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7356_ fd._2446_ fd._2448_ VGND VGND VPWR VPWR fd._2619_ sky130_fd_sc_hd__xnor2_1
XFILLER_257_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4568_ fd._2155_ fd._3661_ VGND VGND VPWR VPWR fd._3662_ sky130_fd_sc_hd__nor2_1
XFILLER_233_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6307_ fd._0846_ fd._1464_ VGND VGND VPWR VPWR fd._1465_ sky130_fd_sc_hd__nand2_1
XFILLER_238_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7287_ fd._2373_ fd._2542_ fd._2505_ VGND VGND VPWR VPWR fd._2543_ sky130_fd_sc_hd__mux2_1
XFILLER_42_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4499_ fd._3590_ VGND VGND VPWR VPWR fd._3593_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_244_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._6238_ fd._1349_ fd._1387_ fd._1388_ VGND VGND VPWR VPWR fd._1389_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6169_ fd._1061_ fd._1312_ fd._1232_ VGND VGND VPWR VPWR fd._1313_ sky130_fd_sc_hd__mux2_1
XFILLER_164_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_257_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_251_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_255_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_250_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_272_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5540_ fd._0618_ fd._0620_ VGND VGND VPWR VPWR fd._0621_ sky130_fd_sc_hd__xor2_1
XFILLER_152_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_258_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5471_ fd._0543_ fd._0544_ VGND VGND VPWR VPWR fd._0545_ sky130_fd_sc_hd__xor2_1
XTAP_7594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7210_ fd._2457_ VGND VGND VPWR VPWR fd._2458_ sky130_fd_sc_hd__clkinv_4
XFILLER_94_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4422_ fd.b\[3\] fd._1880_ VGND VGND VPWR VPWR fd._3516_ sky130_fd_sc_hd__or2_1
XTAP_6871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8190_ net72 fd.mc\[14\] VGND VGND VPWR VPWR fd.c\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_267_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7141_ fd._1976_ fd._2376_ fd._2379_ fd._2381_ VGND VGND VPWR VPWR fd._2382_ sky130_fd_sc_hd__o31ai_1
Xfd._4353_ fd._2969_ fd._3024_ fd._3057_ VGND VGND VPWR VPWR fd._3068_ sky130_fd_sc_hd__a21o_1
XFILLER_281_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_282_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7072_ fd._2234_ fd._2305_ fd._2238_ VGND VGND VPWR VPWR fd._2306_ sky130_fd_sc_hd__o21ai_1
Xfd._4284_ fd._2199_ fd._2276_ fd._2265_ VGND VGND VPWR VPWR fd._2309_ sky130_fd_sc_hd__o21ai_1
XFILLER_235_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6023_ fd._0889_ fd._1151_ fd._1047_ VGND VGND VPWR VPWR fd._1152_ sky130_fd_sc_hd__mux2_1
XFILLER_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_280_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_280_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7974_ fd._0504_ fd._3297_ VGND VGND VPWR VPWR fd._3298_ sky130_fd_sc_hd__and2_1
XFILLER_202_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6925_ fd._1966_ fd._1982_ VGND VGND VPWR VPWR fd._2145_ sky130_fd_sc_hd__nor2_1
XFILLER_148_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6856_ fd._1330_ fd._1894_ VGND VGND VPWR VPWR fd._2069_ sky130_fd_sc_hd__and2_1
XFILLER_11_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5807_ fd._0089_ fd._0914_ VGND VGND VPWR VPWR fd._0915_ sky130_fd_sc_hd__or2_1
XFILLER_116_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6787_ fd._1992_ VGND VGND VPWR VPWR fd._1993_ sky130_fd_sc_hd__inv_2
XFILLER_85_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5738_ fd._0806_ fd._0810_ fd._0838_ VGND VGND VPWR VPWR fd._0839_ sky130_fd_sc_hd__and3_1
XFILLER_103_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_277_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5669_ fd._0482_ fd._0762_ VGND VGND VPWR VPWR fd._0763_ sky130_fd_sc_hd__or2_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7408_ fd._2670_ fd._2675_ VGND VGND VPWR VPWR fd._2676_ sky130_fd_sc_hd__nand2_4
XTAP_4209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7339_ fd._1872_ fd._2598_ VGND VGND VPWR VPWR fd._2600_ sky130_fd_sc_hd__and2_1
XFILLER_84_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_279_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_279_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_257_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_249_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_264_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_262_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4971_ fd._3827_ fd._4066_ fd._3960_ VGND VGND VPWR VPWR fd._4067_ sky130_fd_sc_hd__mux2_1
XFILLER_223_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._6710_ fd._1848_ fd._1905_ fd._1907_ VGND VGND VPWR VPWR fd._1908_ sky130_fd_sc_hd__a21oi_2
XFILLER_145_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_258_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7690_ fd._2899_ fd._2985_ VGND VGND VPWR VPWR fd._2986_ sky130_fd_sc_hd__nand2_1
XFILLER_32_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6641_ fd._1831_ fd._1820_ VGND VGND VPWR VPWR fd._1832_ sky130_fd_sc_hd__nor2_1
XFILLER_67_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6572_ fd._1751_ fd._1755_ VGND VGND VPWR VPWR fd._1756_ sky130_fd_sc_hd__and2_1
XFILLER_154_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5523_ fd._0470_ fd._0396_ VGND VGND VPWR VPWR fd._0602_ sky130_fd_sc_hd__or2b_1
XFILLER_140_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8242_ net74 net23 VGND VGND VPWR VPWR fd.b\[2\] sky130_fd_sc_hd__dfxtp_2
XFILLER_234_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5454_ fd._3708_ VGND VGND VPWR VPWR fd._0526_ sky130_fd_sc_hd__buf_6
XFILLER_132_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_1436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4405_ fd._1759_ fd._2056_ VGND VGND VPWR VPWR fd._3499_ sky130_fd_sc_hd__nand2_1
XFILLER_228_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8173_ fd._3485_ fd._3486_ VGND VGND VPWR VPWR fd._3487_ sky130_fd_sc_hd__xnor2_1
XFILLER_66_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5385_ fd._0279_ fd._0449_ VGND VGND VPWR VPWR fd._0451_ sky130_fd_sc_hd__xor2_1
XFILLER_110_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_269_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7124_ fd._2174_ fd._2362_ VGND VGND VPWR VPWR fd._2363_ sky130_fd_sc_hd__nor2_1
XFILLER_66_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4336_ fd._2815_ fd._2870_ fd._1231_ VGND VGND VPWR VPWR fd._2881_ sky130_fd_sc_hd__mux2_1
XFILLER_48_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_282_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_270_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7055_ fd._1685_ fd._2286_ VGND VGND VPWR VPWR fd._2288_ sky130_fd_sc_hd__nor2_1
Xfd._4267_ fd._0428_ fd._2111_ VGND VGND VPWR VPWR fd._2122_ sky130_fd_sc_hd__and2_1
XFILLER_35_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6006_ fd._0897_ fd._0953_ fd._0959_ VGND VGND VPWR VPWR fd._1134_ sky130_fd_sc_hd__and3_1
XFILLER_165_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4198_ fd._0835_ fd._0956_ VGND VGND VPWR VPWR fd._1363_ sky130_fd_sc_hd__and2_1
XFILLER_222_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7957_ fd._3273_ fd._3274_ fd._3275_ fd._3279_ VGND VGND VPWR VPWR fd._3280_ sky130_fd_sc_hd__a31o_1
XFILLER_109_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6908_ fd._2124_ fd._2125_ VGND VGND VPWR VPWR fd._2126_ sky130_fd_sc_hd__nor2_1
XFILLER_135_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7888_ fd._1685_ fd._3095_ VGND VGND VPWR VPWR fd._3204_ sky130_fd_sc_hd__or2_1
XFILLER_190_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6839_ fd._1904_ fd._1852_ fd._1900_ VGND VGND VPWR VPWR fd._2050_ sky130_fd_sc_hd__and3_1
XFILLER_151_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_1527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_277_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_225_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_1667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_1463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_270_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5170_ fd._0213_ fd._0022_ fd._0067_ VGND VGND VPWR VPWR fd._0214_ sky130_fd_sc_hd__mux2_1
XTAP_4573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4121_ fd.b\[11\] fd.a\[11\] VGND VGND VPWR VPWR fd._0516_ sky130_fd_sc_hd__xor2_1
XFILLER_252_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._7811_ fd._3103_ fd._3118_ VGND VGND VPWR VPWR fd._3119_ sky130_fd_sc_hd__and2_1
XFILLER_9_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_277_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4954_ fd._3841_ fd._3916_ VGND VGND VPWR VPWR fd._4048_ sky130_fd_sc_hd__xor2_1
XFILLER_199_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._7742_ fd._2481_ fd._3042_ VGND VGND VPWR VPWR fd._3043_ sky130_fd_sc_hd__xnor2_1
XFILLER_117_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_277_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7673_ fd._2742_ fd._2770_ fd._2737_ VGND VGND VPWR VPWR fd._2967_ sky130_fd_sc_hd__a21oi_1
XFILLER_133_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4885_ fd._3892_ fd._3978_ fd._3959_ VGND VGND VPWR VPWR fd._3979_ sky130_fd_sc_hd__mux2_2
XFILLER_86_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6624_ fd._1720_ VGND VGND VPWR VPWR fd._1813_ sky130_fd_sc_hd__buf_6
XFILLER_138_1634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6555_ fd._1565_ VGND VGND VPWR VPWR fd._1738_ sky130_fd_sc_hd__clkinv_2
XFILLER_141_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_259_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5506_ fd._0967_ fd._0583_ VGND VGND VPWR VPWR fd._0584_ sky130_fd_sc_hd__xnor2_1
XFILLER_141_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_274_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_253_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6486_ fd._1648_ fd._1658_ fd._1661_ VGND VGND VPWR VPWR fd._1662_ sky130_fd_sc_hd__o21ai_2
XFILLER_228_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_268_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8225_ net70 net9 VGND VGND VPWR VPWR fd.a\[17\] sky130_fd_sc_hd__dfxtp_1
Xfd._5437_ fd._0327_ fd._0507_ VGND VGND VPWR VPWR fd._0508_ sky130_fd_sc_hd__and2_1
XFILLER_283_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_269_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8156_ fd._3460_ fd._3464_ fd._3468_ VGND VGND VPWR VPWR fd._3471_ sky130_fd_sc_hd__o21a_1
XFILLER_23_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5368_ fd._0125_ fd._0431_ VGND VGND VPWR VPWR fd._0432_ sky130_fd_sc_hd__nor2_1
XFILLER_67_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_269_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_270_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7107_ fd._1173_ fd._2344_ VGND VGND VPWR VPWR fd._2345_ sky130_fd_sc_hd__nand2_1
XFILLER_110_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4319_ fd.b\[17\] fd._2683_ VGND VGND VPWR VPWR fd._2694_ sky130_fd_sc_hd__and2_1
Xfd._8087_ fd._1423_ fd._1617_ fd._3411_ VGND VGND VPWR VPWR fd._3412_ sky130_fd_sc_hd__mux2_1
XFILLER_39_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_270_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._5299_ fd._3716_ fd._0355_ VGND VGND VPWR VPWR fd._0356_ sky130_fd_sc_hd__or2_1
XFILLER_42_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7038_ fd._2267_ fd._2268_ VGND VGND VPWR VPWR fd._2269_ sky130_fd_sc_hd__nor2_1
XFILLER_51_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_8828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_278_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_271_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_265_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4670_ fd._3035_ fd._3598_ fd._3600_ VGND VGND VPWR VPWR fd._3764_ sky130_fd_sc_hd__o21bai_1
XFILLER_237_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_272_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6340_ fd._0131_ fd._1428_ VGND VGND VPWR VPWR fd._1501_ sky130_fd_sc_hd__nand2_1
XFILLER_123_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6271_ fd._1088_ fd._1424_ VGND VGND VPWR VPWR fd._1425_ sky130_fd_sc_hd__xnor2_1
XFILLER_283_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 io_in[16] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
XTAP_5082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._8010_ fd._3110_ fd._3117_ fd._3202_ fd._3334_ VGND VGND VPWR VPWR fd._3338_ sky130_fd_sc_hd__o22ai_2
XFILLER_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5222_ fd._0231_ fd._0267_ fd._0270_ VGND VGND VPWR VPWR fd._0271_ sky130_fd_sc_hd__mux2_1
XTAP_5093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_280_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5153_ fd._0194_ VGND VGND VPWR VPWR fd._0195_ sky130_fd_sc_hd__inv_2
XFILLER_24_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4104_ fd.b\[2\] fd.a\[2\] VGND VGND VPWR VPWR fd._0329_ sky130_fd_sc_hd__and2b_1
XFILLER_33_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5084_ fd._3869_ fd._0118_ VGND VGND VPWR VPWR fd._0119_ sky130_fd_sc_hd__and2_1
XFILLER_75_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5986_ fd._1104_ fd._1109_ fd._1111_ VGND VGND VPWR VPWR fd._1112_ sky130_fd_sc_hd__o21bai_1
XFILLER_257_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_277_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7725_ fd._3023_ VGND VGND VPWR VPWR fd._3025_ sky130_fd_sc_hd__clkinv_2
Xfd._4937_ fd._4030_ fd._3894_ VGND VGND VPWR VPWR fd._4031_ sky130_fd_sc_hd__xnor2_1
XFILLER_118_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_255_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4868_ fd._3789_ fd._3941_ fd._3961_ VGND VGND VPWR VPWR fd._3962_ sky130_fd_sc_hd__mux2_1
Xfd._7656_ fd._2948_ fd._2764_ VGND VGND VPWR VPWR fd._2949_ sky130_fd_sc_hd__nor2_1
XFILLER_273_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_255_1644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_251_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6607_ fd._0343_ fd._1793_ VGND VGND VPWR VPWR fd._1795_ sky130_fd_sc_hd__nor2_1
XFILLER_138_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_255_1688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._4799_ fd._3708_ fd._3892_ VGND VGND VPWR VPWR fd._3893_ sky130_fd_sc_hd__nor2_1
XFILLER_138_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._7587_ fd._2871_ fd._2872_ fd._2856_ fd._2864_ VGND VGND VPWR VPWR fd._2873_ sky130_fd_sc_hd__a22o_1
XFILLER_141_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6538_ fd._1626_ fd._1644_ fd._1718_ VGND VGND VPWR VPWR fd._1719_ sky130_fd_sc_hd__nand3_4
XFILLER_25_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6469_ fd._1165_ fd._1630_ VGND VGND VPWR VPWR fd._1643_ sky130_fd_sc_hd__nor2_1
XFILLER_74_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8208_ net74 net1 VGND VGND VPWR VPWR fd.a\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_28_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_283_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_284_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8139_ fd._3440_ fd._3445_ fd._3452_ VGND VGND VPWR VPWR fd._3454_ sky130_fd_sc_hd__o21a_1
XFILLER_215_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_282_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_273_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_1546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5840_ fd._0950_ VGND VGND VPWR VPWR fd._0951_ sky130_fd_sc_hd__inv_2
XFILLER_278_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_259_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5771_ fd._0653_ fd._0749_ fd._0754_ VGND VGND VPWR VPWR fd._0875_ sky130_fd_sc_hd__nand3_1
XFILLER_278_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4722_ fd._3815_ fd._3740_ fd._3788_ VGND VGND VPWR VPWR fd._3816_ sky130_fd_sc_hd__mux2_1
XFILLER_155_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7510_ fd._2517_ fd._2523_ fd._2565_ fd._2515_ VGND VGND VPWR VPWR fd._2788_ sky130_fd_sc_hd__a31o_1
XFILLER_13_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4653_ fd._3637_ fd._3746_ VGND VGND VPWR VPWR fd._3747_ sky130_fd_sc_hd__nand2_1
XFILLER_174_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7441_ fd._2710_ fd._2711_ VGND VGND VPWR VPWR fd._2712_ sky130_fd_sc_hd__nor2_1
XFILLER_29_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7372_ fd._2481_ fd._2635_ VGND VGND VPWR VPWR fd._2636_ sky130_fd_sc_hd__nand2_1
XFILLER_135_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4584_ fd._3676_ fd._3677_ VGND VGND VPWR VPWR fd._3678_ sky130_fd_sc_hd__xnor2_1
XFILLER_284_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6323_ fd._4055_ fd._1477_ fd._1481_ VGND VGND VPWR VPWR fd._1482_ sky130_fd_sc_hd__mux2_1
XFILLER_110_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_1372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6254_ fd._1189_ fd._1216_ VGND VGND VPWR VPWR fd._1406_ sky130_fd_sc_hd__nand2_1
XFILLER_2_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5205_ fd._3689_ fd._0061_ fd._0062_ fd._0235_ fd._0239_ VGND VGND VPWR VPWR fd._0253_
+ sky130_fd_sc_hd__a221o_1
XFILLER_38_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6185_ fd._1309_ fd._1078_ VGND VGND VPWR VPWR fd._1331_ sky130_fd_sc_hd__xor2_1
XFILLER_64_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_1408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5136_ fd._0168_ fd._0173_ fd._0176_ VGND VGND VPWR VPWR fd._0177_ sky130_fd_sc_hd__a21o_1
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5067_ fd._3999_ fd._4015_ VGND VGND VPWR VPWR fd._0101_ sky130_fd_sc_hd__nand2_1
XFILLER_221_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_13 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5969_ fd._0916_ fd._1082_ VGND VGND VPWR VPWR fd._1093_ sky130_fd_sc_hd__or2_1
XFILLER_273_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7708_ fd._0382_ fd._3005_ VGND VGND VPWR VPWR fd._3006_ sky130_fd_sc_hd__or2_1
XFILLER_31_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7639_ fd._2748_ VGND VGND VPWR VPWR fd._2930_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_47_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xuser_project_wrapper_190 VGND VGND VPWR VPWR user_project_wrapper_190/HI la_data_out[68]
+ sky130_fd_sc_hd__conb_1
XFILLER_62_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_251_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_276_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_271_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_9145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_1506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_278_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_266_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_281_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7990_ fd._3315_ fd._3186_ VGND VGND VPWR VPWR fd._3316_ sky130_fd_sc_hd__xnor2_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6941_ fd._1966_ fd._2161_ VGND VGND VPWR VPWR fd._2162_ sky130_fd_sc_hd__nor2_1
XFILLER_72_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1690 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput11 io_in[19] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_2
XFILLER_238_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6872_ fd._2085_ fd._1882_ VGND VGND VPWR VPWR fd._2086_ sky130_fd_sc_hd__xnor2_1
XFILLER_141_1652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput22 io_in[29] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
XFILLER_141_1663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput33 wb_clk_i VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_16
Xfd._5823_ fd._0910_ fd._0931_ VGND VGND VPWR VPWR fd._0932_ sky130_fd_sc_hd__nand2_1
XFILLER_162_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5754_ fd._0786_ fd._0855_ VGND VGND VPWR VPWR fd._0856_ sky130_fd_sc_hd__or2_1
XFILLER_192_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4705_ fd._3796_ fd._3797_ VGND VGND VPWR VPWR fd._3799_ sky130_fd_sc_hd__nand2_1
Xfd._5685_ fd._0755_ fd._0756_ fd._0763_ fd._0778_ fd._0779_ VGND VGND VPWR VPWR fd._0781_
+ sky130_fd_sc_hd__a311oi_4
XFILLER_192_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7424_ fd._1666_ fd._2604_ VGND VGND VPWR VPWR fd._2693_ sky130_fd_sc_hd__nand2_1
XFILLER_44_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4636_ fd._3416_ fd._3729_ fd._3625_ VGND VGND VPWR VPWR fd._3730_ sky130_fd_sc_hd__mux2_1
XFILLER_269_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_284_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4567_ fd._3502_ fd._3660_ fd._3624_ VGND VGND VPWR VPWR fd._3661_ sky130_fd_sc_hd__mux2_1
XFILLER_229_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7355_ fd._2443_ VGND VGND VPWR VPWR fd._2618_ sky130_fd_sc_hd__clkinv_2
XFILLER_57_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6306_ fd._1460_ fd._1463_ fd._1422_ VGND VGND VPWR VPWR fd._1464_ sky130_fd_sc_hd__mux2_1
XFILLER_96_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_285_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_226_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7286_ fd._2539_ fd._2541_ VGND VGND VPWR VPWR fd._2542_ sky130_fd_sc_hd__xor2_1
XFILLER_2_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._4498_ fd._3577_ fd._3582_ fd._3590_ fd._3591_ VGND VGND VPWR VPWR fd._3592_ sky130_fd_sc_hd__o31a_1
XFILLER_211_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6237_ fd._1210_ fd._1340_ fd._1348_ VGND VGND VPWR VPWR fd._1388_ sky130_fd_sc_hd__and3_1
XFILLER_246_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_253_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6168_ fd._1310_ fd._1311_ VGND VGND VPWR VPWR fd._1312_ sky130_fd_sc_hd__xnor2_1
XFILLER_164_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5119_ fd._3982_ fd._4028_ fd._0157_ VGND VGND VPWR VPWR fd._0158_ sky130_fd_sc_hd__and3_1
XFILLER_0_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6099_ fd._1137_ fd._1235_ fd._1223_ VGND VGND VPWR VPWR fd._1236_ sky130_fd_sc_hd__mux2_1
XFILLER_146_1552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_264_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_262_1286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_275_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_256_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5470_ fd._0349_ fd._0348_ VGND VGND VPWR VPWR fd._0544_ sky130_fd_sc_hd__or2b_1
XFILLER_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4421_ fd._1935_ fd._2001_ VGND VGND VPWR VPWR fd._3515_ sky130_fd_sc_hd__and2_1
XTAP_6861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7140_ fd._1970_ fd._2250_ fd._2321_ fd._2377_ VGND VGND VPWR VPWR fd._2381_ sky130_fd_sc_hd__a31o_1
XFILLER_282_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4352_ fd._2892_ fd._3046_ VGND VGND VPWR VPWR fd._3057_ sky130_fd_sc_hd__nand2_1
XFILLER_212_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_282_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7071_ fd._2233_ fd._2109_ VGND VGND VPWR VPWR fd._2305_ sky130_fd_sc_hd__nor2_1
XFILLER_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4283_ fd._2265_ fd._2287_ VGND VGND VPWR VPWR fd._2298_ sky130_fd_sc_hd__nand2_1
XFILLER_235_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_281_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6022_ fd._1149_ fd._1150_ VGND VGND VPWR VPWR fd._1151_ sky130_fd_sc_hd__xnor2_1
XFILLER_267_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_280_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7973_ fd._3151_ fd._3296_ fd._3239_ VGND VGND VPWR VPWR fd._3297_ sky130_fd_sc_hd__mux2_1
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_280_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6924_ fd._2142_ fd._1955_ VGND VGND VPWR VPWR fd._2143_ sky130_fd_sc_hd__or2_1
XFILLER_147_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6855_ fd._1864_ fd._1892_ VGND VGND VPWR VPWR fd._2068_ sky130_fd_sc_hd__or2_1
XFILLER_163_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5806_ fd._0665_ fd._0913_ fd._0801_ VGND VGND VPWR VPWR fd._0914_ sky130_fd_sc_hd__mux2_1
XFILLER_162_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._6786_ fd._1932_ fd._1925_ VGND VGND VPWR VPWR fd._1992_ sky130_fd_sc_hd__and2b_1
XFILLER_116_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5737_ fd._0819_ fd._0836_ fd._0837_ fd._0817_ VGND VGND VPWR VPWR fd._0838_ sky130_fd_sc_hd__a211o_1
XFILLER_171_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5668_ fd._0760_ fd._0761_ fd._0672_ fd._0757_ VGND VGND VPWR VPWR fd._0762_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_135_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7407_ fd._1816_ fd._2665_ fd._2667_ fd._2674_ VGND VGND VPWR VPWR fd._2675_ sky130_fd_sc_hd__o31a_4
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_281_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4619_ fd._3469_ fd._3653_ VGND VGND VPWR VPWR fd._3713_ sky130_fd_sc_hd__nand2_1
XFILLER_258_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5599_ fd._0526_ fd._0675_ VGND VGND VPWR VPWR fd._0686_ sky130_fd_sc_hd__nor2_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._7338_ fd._1872_ fd._2598_ VGND VGND VPWR VPWR fd._2599_ sky130_fd_sc_hd__or2_1
XFILLER_6_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7269_ fd._1219_ fd._2522_ VGND VGND VPWR VPWR fd._2523_ sky130_fd_sc_hd__nand2_1
XFILLER_2_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_260_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_246_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_279_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_264_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_263_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_281_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4970_ fd._4065_ VGND VGND VPWR VPWR fd._4066_ sky130_fd_sc_hd__clkinv_2
XFILLER_33_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6640_ fd._2738_ fd._1830_ VGND VGND VPWR VPWR fd._1831_ sky130_fd_sc_hd__nor2_1
XFILLER_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._6571_ fd._1581_ fd._1754_ fd._1719_ VGND VGND VPWR VPWR fd._1755_ sky130_fd_sc_hd__mux2_1
XFILLER_10_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_275_1499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5522_ fd._0482_ fd._0600_ VGND VGND VPWR VPWR fd._0601_ sky130_fd_sc_hd__nor2_1
XFILLER_49_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8241_ net74 net12 VGND VGND VPWR VPWR fd.b\[1\] sky130_fd_sc_hd__dfxtp_4
XTAP_7392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5453_ fd._0514_ fd._0521_ fd._0524_ fd._0512_ VGND VGND VPWR VPWR fd._0525_ sky130_fd_sc_hd__a31oi_2
XFILLER_79_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4404_ fd._3490_ fd._3496_ fd._3497_ VGND VGND VPWR VPWR fd._3498_ sky130_fd_sc_hd__a21o_1
XFILLER_171_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5384_ fd._0420_ fd._0413_ fd._0416_ VGND VGND VPWR VPWR fd._0449_ sky130_fd_sc_hd__o21ai_1
Xfd._8172_ fd._3478_ fd._3481_ fd._3476_ VGND VGND VPWR VPWR fd._3486_ sky130_fd_sc_hd__o21a_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4335_ fd._1011_ fd._2859_ VGND VGND VPWR VPWR fd._2870_ sky130_fd_sc_hd__xnor2_1
XFILLER_243_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7123_ fd._1958_ fd._2173_ VGND VGND VPWR VPWR fd._2362_ sky130_fd_sc_hd__nor2_1
XFILLER_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_242_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4266_ fd._0483_ fd._2100_ fd._1209_ VGND VGND VPWR VPWR fd._2111_ sky130_fd_sc_hd__mux2_1
XFILLER_169_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7054_ fd._2270_ fd._2275_ fd._2285_ fd._2277_ VGND VGND VPWR VPWR fd._2286_ sky130_fd_sc_hd__a211oi_1
XFILLER_165_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_251_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6005_ fd._0726_ fd._1127_ fd._1131_ VGND VGND VPWR VPWR fd._1133_ sky130_fd_sc_hd__mux2_1
XFILLER_23_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4197_ fd.b\[19\] VGND VGND VPWR VPWR fd._1352_ sky130_fd_sc_hd__buf_6
XFILLER_165_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_280_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7956_ fd._3240_ fd._3278_ VGND VGND VPWR VPWR fd._3279_ sky130_fd_sc_hd__nand2_1
XFILLER_17_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6907_ fd._1872_ fd._2123_ VGND VGND VPWR VPWR fd._2125_ sky130_fd_sc_hd__nor2_1
XFILLER_108_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7887_ fd._3127_ fd._3197_ fd._3202_ fd._3121_ VGND VGND VPWR VPWR fd._3203_ sky130_fd_sc_hd__a211o_1
XFILLER_11_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._6838_ fd._1852_ fd._1900_ fd._1904_ VGND VGND VPWR VPWR fd._2049_ sky130_fd_sc_hd__a21oi_1
XFILLER_190_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6769_ fd._1961_ fd._1972_ VGND VGND VPWR VPWR fd._1973_ sky130_fd_sc_hd__and2b_1
XFILLER_143_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_269_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_249_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4120_ fd._0428_ fd._0439_ fd._0208_ fd._0472_ fd._0494_ VGND VGND VPWR VPWR fd._0505_
+ sky130_fd_sc_hd__o221a_1
XFILLER_251_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7810_ fd._2076_ fd._3102_ VGND VGND VPWR VPWR fd._3118_ sky130_fd_sc_hd__nand2_1
XFILLER_14_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7741_ fd._2828_ fd._3041_ fd._2877_ VGND VGND VPWR VPWR fd._3042_ sky130_fd_sc_hd__mux2_1
Xfd._4953_ fd._4042_ fd._3833_ fd._4046_ VGND VGND VPWR VPWR fd._4047_ sky130_fd_sc_hd__mux2_1
XFILLER_146_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7672_ fd._2737_ fd._2742_ fd._2770_ VGND VGND VPWR VPWR fd._2966_ sky130_fd_sc_hd__and3_1
Xfd._4884_ fd._3888_ fd._3977_ VGND VGND VPWR VPWR fd._3978_ sky130_fd_sc_hd__xnor2_1
XFILLER_12_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6623_ fd._1807_ fd._1641_ VGND VGND VPWR VPWR fd._1812_ sky130_fd_sc_hd__xnor2_1
XFILLER_132_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6554_ fd._0928_ fd._1735_ VGND VGND VPWR VPWR fd._1736_ sky130_fd_sc_hd__nor2_1
XFILLER_119_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_262_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_259_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5505_ fd._0383_ fd._0581_ fd._0452_ VGND VGND VPWR VPWR fd._0583_ sky130_fd_sc_hd__mux2_1
XFILLER_119_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6485_ fd._1451_ VGND VGND VPWR VPWR fd._1661_ sky130_fd_sc_hd__buf_6
XFILLER_136_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8224_ net71 net8 VGND VGND VPWR VPWR fd.a\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_269_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5436_ fd._0324_ fd._0325_ VGND VGND VPWR VPWR fd._0507_ sky130_fd_sc_hd__or2_1
XFILLER_210_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_267_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_269_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8155_ fd._3460_ fd._3464_ fd._3468_ VGND VGND VPWR VPWR fd._3470_ sky130_fd_sc_hd__nor3_1
XFILLER_82_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5367_ fd._0253_ fd._0255_ VGND VGND VPWR VPWR fd._0431_ sky130_fd_sc_hd__nand2_1
XFILLER_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_283_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_270_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_269_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7106_ fd._2139_ fd._2343_ fd._2322_ VGND VGND VPWR VPWR fd._2344_ sky130_fd_sc_hd__mux2_1
Xfd._4318_ fd._0043_ fd._1374_ fd._1231_ VGND VGND VPWR VPWR fd._2683_ sky130_fd_sc_hd__mux2_1
XFILLER_82_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8086_ fd._3189_ VGND VGND VPWR VPWR fd._3411_ sky130_fd_sc_hd__buf_4
Xfd._5298_ fd._0152_ fd._0354_ fd._0269_ VGND VGND VPWR VPWR fd._0355_ sky130_fd_sc_hd__mux2_1
XFILLER_93_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7037_ fd._2076_ fd._2266_ VGND VGND VPWR VPWR fd._2268_ sky130_fd_sc_hd__nor2_1
XFILLER_35_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4249_ fd._1902_ fd._1913_ fd._1209_ VGND VGND VPWR VPWR fd._1924_ sky130_fd_sc_hd__mux2_1
XFILLER_184_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_1663 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_260_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7939_ fd._3257_ fd._3259_ VGND VGND VPWR VPWR fd._3260_ sky130_fd_sc_hd__xnor2_1
XFILLER_17_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_276_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_1601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_261_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_1523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_257_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6270_ fd._1306_ fd._1421_ fd._1423_ VGND VGND VPWR VPWR fd._1424_ sky130_fd_sc_hd__mux2_1
XTAP_5050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput9 io_in[17] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
Xfd._5221_ fd._0269_ VGND VGND VPWR VPWR fd._0270_ sky130_fd_sc_hd__buf_6
XTAP_5083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5152_ fd._0191_ fd._0192_ fd._0067_ fd._0193_ VGND VGND VPWR VPWR fd._0194_ sky130_fd_sc_hd__o31a_1
XFILLER_248_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_1663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4103_ fd._0296_ VGND VGND VPWR VPWR fd._0318_ sky130_fd_sc_hd__buf_4
XFILLER_205_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5083_ fd._0117_ fd._0114_ fd._0059_ VGND VGND VPWR VPWR fd._0118_ sky130_fd_sc_hd__mux2_1
XFILLER_209_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_233_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5985_ fd._0541_ fd._1108_ VGND VGND VPWR VPWR fd._1111_ sky130_fd_sc_hd__and2_1
XFILLER_277_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7724_ fd._3022_ fd._2865_ VGND VGND VPWR VPWR fd._3023_ sky130_fd_sc_hd__xnor2_1
Xfd._4936_ fd._3897_ fd._3973_ fd._3851_ VGND VGND VPWR VPWR fd._4030_ sky130_fd_sc_hd__o21a_1
XFILLER_238_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_1571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7655_ fd._2763_ fd._2945_ VGND VGND VPWR VPWR fd._2948_ sky130_fd_sc_hd__nor2_1
XFILLER_133_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4867_ fd._3960_ VGND VGND VPWR VPWR fd._3961_ sky130_fd_sc_hd__buf_6
XFILLER_173_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6606_ fd._0343_ fd._1793_ VGND VGND VPWR VPWR fd._1794_ sky130_fd_sc_hd__nand2_1
XFILLER_114_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_1629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._7586_ fd._2674_ fd._2869_ fd._2665_ VGND VGND VPWR VPWR fd._2872_ sky130_fd_sc_hd__o21ai_1
XFILLER_86_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4798_ fd._3889_ fd._3800_ fd._3890_ fd._3891_ VGND VGND VPWR VPWR fd._3892_ sky130_fd_sc_hd__a31oi_2
XFILLER_87_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6537_ fd._1703_ fd._1709_ fd._1712_ fd._1713_ fd._1717_ VGND VGND VPWR VPWR fd._1718_
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_141_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._6468_ fd._1618_ fd._1641_ VGND VGND VPWR VPWR fd._1642_ sky130_fd_sc_hd__nand2_1
XFILLER_228_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8207_ net69 fd.sc VGND VGND VPWR VPWR fd.c\[31\] sky130_fd_sc_hd__dfxtp_1
Xfd._5419_ fd._0484_ fd._0487_ fd._0452_ VGND VGND VPWR VPWR fd._0488_ sky130_fd_sc_hd__mux2_1
XFILLER_67_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6399_ fd._1559_ fd._1565_ VGND VGND VPWR VPWR fd._1566_ sky130_fd_sc_hd__nand2_1
XFILLER_215_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8138_ fd._3440_ fd._3445_ fd._3452_ VGND VGND VPWR VPWR fd._3453_ sky130_fd_sc_hd__nor3_1
XFILLER_83_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_270_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._8069_ fd._3400_ VGND VGND VPWR VPWR fd.mc\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_97_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_223_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_260_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_260_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_279_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_278_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_281_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_259_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5770_ fd._0861_ fd._0870_ fd._0873_ VGND VGND VPWR VPWR fd._0874_ sky130_fd_sc_hd__nand3_2
XFILLER_41_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_278_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4721_ fd._3738_ fd._3814_ VGND VGND VPWR VPWR fd._3815_ sky130_fd_sc_hd__xnor2_1
XFILLER_170_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_276_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7440_ fd._1797_ fd._2709_ VGND VGND VPWR VPWR fd._2711_ sky130_fd_sc_hd__nor2_1
Xfd._4652_ fd._1253_ fd._3636_ VGND VGND VPWR VPWR fd._3746_ sky130_fd_sc_hd__nand2_1
XFILLER_237_1364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7371_ fd._2425_ fd._2634_ fd._2623_ VGND VGND VPWR VPWR fd._2635_ sky130_fd_sc_hd__mux2_1
XFILLER_257_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4583_ fd._3531_ fd._3540_ VGND VGND VPWR VPWR fd._3677_ sky130_fd_sc_hd__or2b_1
XFILLER_2_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6322_ fd._1478_ fd._1480_ VGND VGND VPWR VPWR fd._1481_ sky130_fd_sc_hd__xnor2_1
XFILLER_96_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_250_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_250_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6253_ fd._1371_ fd._1377_ fd._1404_ fd._1369_ VGND VGND VPWR VPWR fd._1405_ sky130_fd_sc_hd__a31o_1
XFILLER_133_1384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5204_ fd._0240_ fd._0250_ VGND VGND VPWR VPWR fd._0251_ sky130_fd_sc_hd__and2_1
XFILLER_20_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_266_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6184_ fd._1327_ fd._1328_ VGND VGND VPWR VPWR fd._1329_ sky130_fd_sc_hd__nor2_1
XTAP_4190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_252_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5135_ fd._0758_ fd._0174_ VGND VGND VPWR VPWR fd._0176_ sky130_fd_sc_hd__nor2_1
XFILLER_94_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5066_ fd._0097_ fd._0099_ VGND VGND VPWR VPWR fd._0100_ sky130_fd_sc_hd__nor2_1
XFILLER_127_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_14 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5968_ fd._1087_ fd._1091_ VGND VGND VPWR VPWR fd._1092_ sky130_fd_sc_hd__or2_1
XFILLER_179_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7707_ fd._2697_ fd._3004_ fd._2875_ VGND VGND VPWR VPWR fd._3005_ sky130_fd_sc_hd__mux2_1
Xfd._4919_ fd._3688_ fd._4006_ fd._4009_ fd._4012_ VGND VGND VPWR VPWR fd._4013_ sky130_fd_sc_hd__o31a_1
XFILLER_118_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5899_ fd._0638_ fd._0830_ VGND VGND VPWR VPWR fd._1016_ sky130_fd_sc_hd__nor2_1
XFILLER_133_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7638_ fd._2927_ fd._2928_ VGND VGND VPWR VPWR fd._2929_ sky130_fd_sc_hd__nor2_1
XTAP_6509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_project_wrapper_180 VGND VGND VPWR VPWR user_project_wrapper_180/HI la_data_out[58]
+ sky130_fd_sc_hd__conb_1
XFILLER_216_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_project_wrapper_191 VGND VGND VPWR VPWR user_project_wrapper_191/HI la_data_out[69]
+ sky130_fd_sc_hd__conb_1
XFILLER_47_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7569_ fd._2852_ fd._2668_ VGND VGND VPWR VPWR fd._2853_ sky130_fd_sc_hd__nand2_1
XFILLER_142_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_276_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_275_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_263_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_255_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_9135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_8445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_279_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_281_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_1600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_1442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6940_ fd._1958_ fd._1965_ VGND VGND VPWR VPWR fd._2161_ sky130_fd_sc_hd__nor2_1
XFILLER_124_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6871_ fd._1796_ fd._1799_ fd._1883_ VGND VGND VPWR VPWR fd._2085_ sky130_fd_sc_hd__o21a_1
XFILLER_198_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput12 io_in[1] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_4
XFILLER_30_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput23 io_in[2] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_4
Xfd._5822_ fd._0662_ fd._0908_ VGND VGND VPWR VPWR fd._0931_ sky130_fd_sc_hd__nand2_1
XFILLER_141_1686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5753_ fd._0774_ fd._0854_ fd._0848_ VGND VGND VPWR VPWR fd._0855_ sky130_fd_sc_hd__mux2_1
XFILLER_171_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4704_ fd._3796_ fd._3797_ VGND VGND VPWR VPWR fd._3798_ sky130_fd_sc_hd__or2_1
XFILLER_196_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5684_ fd._0482_ fd._0762_ VGND VGND VPWR VPWR fd._0779_ sky130_fd_sc_hd__and2_1
XFILLER_170_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_1626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7423_ fd._0382_ fd._2691_ VGND VGND VPWR VPWR fd._2692_ sky130_fd_sc_hd__nand2_1
XFILLER_48_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4635_ fd._3638_ fd._3639_ VGND VGND VPWR VPWR fd._3729_ sky130_fd_sc_hd__xnor2_1
XFILLER_139_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_272_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_258_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7354_ fd._2509_ fd._2614_ fd._2615_ VGND VGND VPWR VPWR fd._2616_ sky130_fd_sc_hd__a21o_1
XFILLER_257_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4566_ fd._3657_ fd._3659_ VGND VGND VPWR VPWR fd._3660_ sky130_fd_sc_hd__xnor2_1
XFILLER_284_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6305_ fd._1258_ fd._1461_ VGND VGND VPWR VPWR fd._1463_ sky130_fd_sc_hd__xnor2_1
XFILLER_284_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7285_ fd._1958_ fd._2373_ VGND VGND VPWR VPWR fd._2541_ sky130_fd_sc_hd__xnor2_1
XFILLER_266_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4497_ fd._3589_ fd._3579_ fd._3588_ VGND VGND VPWR VPWR fd._3591_ sky130_fd_sc_hd__a21bo_1
XFILLER_203_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6236_ fd._1384_ fd._1386_ VGND VGND VPWR VPWR fd._1387_ sky130_fd_sc_hd__xnor2_1
XFILLER_26_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_281_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_285_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_253_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6167_ fd._1075_ fd._1062_ VGND VGND VPWR VPWR fd._1311_ sky130_fd_sc_hd__nor2_1
XFILLER_20_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5118_ fd._4034_ fd._4033_ VGND VGND VPWR VPWR fd._0157_ sky130_fd_sc_hd__or2b_1
XFILLER_34_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6098_ fd._1133_ fd._1234_ VGND VGND VPWR VPWR fd._1235_ sky130_fd_sc_hd__xor2_1
XFILLER_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5049_ fd._4027_ fd._0080_ VGND VGND VPWR VPWR fd._0081_ sky130_fd_sc_hd__xnor2_1
XFILLER_221_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_1644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_249_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_268_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_240_1552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4420_ fd._3513_ VGND VGND VPWR VPWR fd._3514_ sky130_fd_sc_hd__inv_2
XTAP_7596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4351_ fd._3035_ fd._2881_ VGND VGND VPWR VPWR fd._3046_ sky130_fd_sc_hd__nand2_1
XFILLER_266_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7070_ fd._2302_ fd._2303_ VGND VGND VPWR VPWR fd._2304_ sky130_fd_sc_hd__nor2_1
XFILLER_130_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._4282_ fd._2276_ VGND VGND VPWR VPWR fd._2287_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_263_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6021_ fd._0891_ fd._0966_ VGND VGND VPWR VPWR fd._1150_ sky130_fd_sc_hd__nand2_1
XFILLER_250_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_250_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_280_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7972_ fd._3294_ fd._3295_ VGND VGND VPWR VPWR fd._3296_ sky130_fd_sc_hd__xnor2_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6923_ fd._0450_ VGND VGND VPWR VPWR fd._2142_ sky130_fd_sc_hd__buf_6
XFILLER_124_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6854_ fd._1275_ fd._2065_ VGND VGND VPWR VPWR fd._2066_ sky130_fd_sc_hd__nor2_1
XFILLER_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_278_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5805_ fd._0668_ fd._0911_ VGND VGND VPWR VPWR fd._0913_ sky130_fd_sc_hd__xnor2_1
XFILLER_116_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6785_ fd._0928_ fd._1989_ VGND VGND VPWR VPWR fd._1991_ sky130_fd_sc_hd__nand2_1
XFILLER_239_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5736_ fd._0807_ fd._0809_ VGND VGND VPWR VPWR fd._0837_ sky130_fd_sc_hd__nor2_1
XFILLER_239_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_1570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_217_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_258_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5667_ fd._0592_ fd._0759_ fd._0672_ VGND VGND VPWR VPWR fd._0761_ sky130_fd_sc_hd__o21a_1
XFILLER_48_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7406_ fd._2472_ fd._2671_ fd._2673_ VGND VGND VPWR VPWR fd._2674_ sky130_fd_sc_hd__o21ai_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_285_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4618_ fd._3651_ fd._3711_ VGND VGND VPWR VPWR fd._3712_ sky130_fd_sc_hd__or2_1
XFILLER_213_1418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5598_ fd._0623_ fd._0630_ fd._0640_ fd._0642_ fd._0645_ VGND VGND VPWR VPWR fd._0685_
+ sky130_fd_sc_hd__a311o_1
XFILLER_57_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7337_ fd._2402_ fd._2597_ fd._2506_ VGND VGND VPWR VPWR fd._2598_ sky130_fd_sc_hd__mux2_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4549_ fd._3430_ fd._3642_ VGND VGND VPWR VPWR fd._3643_ sky130_fd_sc_hd__xor2_1
XFILLER_245_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7268_ fd._2354_ fd._2521_ fd._2505_ VGND VGND VPWR VPWR fd._2522_ sky130_fd_sc_hd__mux2_1
XFILLER_211_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6219_ fd._1362_ fd._1367_ fd._1349_ VGND VGND VPWR VPWR fd._1368_ sky130_fd_sc_hd__mux2_1
XFILLER_285_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_253_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7199_ fd._2444_ fd._2445_ VGND VGND VPWR VPWR fd._2446_ sky130_fd_sc_hd__and2_1
XFILLER_0_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_257_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_270_1523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6570_ fd._1752_ fd._1753_ VGND VGND VPWR VPWR fd._1754_ sky130_fd_sc_hd__xnor2_1
XTAP_8050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5521_ fd._0592_ fd._0594_ fd._0599_ VGND VGND VPWR VPWR fd._0600_ sky130_fd_sc_hd__mux2_1
XFILLER_165_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8240_ net74 net1 VGND VGND VPWR VPWR fd.b\[0\] sky130_fd_sc_hd__dfxtp_2
XTAP_7382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5452_ fd._0430_ fd._0447_ fd._0522_ fd._0523_ VGND VGND VPWR VPWR fd._0524_ sky130_fd_sc_hd__a211o_1
XFILLER_45_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4403_ fd.b\[9\] fd._3489_ VGND VGND VPWR VPWR fd._3497_ sky130_fd_sc_hd__and2_1
XFILLER_234_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_282_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._8171_ fd.b\[30\] fd.a\[30\] VGND VGND VPWR VPWR fd._3485_ sky130_fd_sc_hd__xor2_1
XFILLER_227_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5383_ fd._0430_ fd._0447_ VGND VGND VPWR VPWR fd._0448_ sky130_fd_sc_hd__xnor2_1
XFILLER_39_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7122_ fd._2184_ fd._2187_ VGND VGND VPWR VPWR fd._2361_ sky130_fd_sc_hd__nand2_1
XFILLER_48_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4334_ fd._1055_ fd._2848_ fd._1044_ VGND VGND VPWR VPWR fd._2859_ sky130_fd_sc_hd__a21oi_1
XFILLER_94_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_1503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7053_ fd._2283_ VGND VGND VPWR VPWR fd._2285_ sky130_fd_sc_hd__clkinvlp_2
Xfd._4265_ fd._0186_ fd._2089_ VGND VGND VPWR VPWR fd._2100_ sky130_fd_sc_hd__xnor2_1
XFILLER_251_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6004_ fd._1128_ fd._1130_ VGND VGND VPWR VPWR fd._1131_ sky130_fd_sc_hd__xnor2_2
XFILLER_165_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_251_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4196_ fd.b\[6\] VGND VGND VPWR VPWR fd._1341_ sky130_fd_sc_hd__inv_2
XFILLER_222_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_280_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7955_ fd._3273_ fd._3276_ fd._2751_ VGND VGND VPWR VPWR fd._3278_ sky130_fd_sc_hd__o21ai_1
XFILLER_31_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1580 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6906_ fd._1872_ fd._2123_ VGND VGND VPWR VPWR fd._2124_ sky130_fd_sc_hd__and2_1
XFILLER_163_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7886_ fd._3199_ fd._3201_ VGND VGND VPWR VPWR fd._3202_ sky130_fd_sc_hd__nand2_1
XFILLER_50_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_276_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6837_ fd._2044_ fd._2047_ VGND VGND VPWR VPWR fd._2048_ sky130_fd_sc_hd__nor2_1
XFILLER_117_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_278_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6768_ fd._1585_ fd._1771_ VGND VGND VPWR VPWR fd._1972_ sky130_fd_sc_hd__nand2_1
XFILLER_116_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5719_ fd._0427_ fd._0816_ VGND VGND VPWR VPWR fd._0818_ sky130_fd_sc_hd__and2_1
XFILLER_277_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6699_ fd._1319_ fd._1894_ VGND VGND VPWR VPWR fd._1896_ sky130_fd_sc_hd__nand2_1
XFILLER_154_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_258_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_252_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_265_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_246_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_257_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_249_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_264_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_277_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_249_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7740_ fd._3028_ fd._3040_ VGND VGND VPWR VPWR fd._3041_ sky130_fd_sc_hd__xor2_1
Xfd._4952_ fd._1451_ fd._4045_ VGND VGND VPWR VPWR fd._4046_ sky130_fd_sc_hd__xnor2_1
XFILLER_201_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7671_ fd._2929_ fd._2934_ fd._2964_ fd._2927_ VGND VGND VPWR VPWR fd._2965_ sky130_fd_sc_hd__a31oi_2
Xfd._4883_ fd._3976_ fd._3893_ VGND VGND VPWR VPWR fd._3977_ sky130_fd_sc_hd__nor2_1
XFILLER_199_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6622_ fd._1625_ fd._1809_ fd._1618_ VGND VGND VPWR VPWR fd._1811_ sky130_fd_sc_hd__a21o_1
XFILLER_154_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6553_ fd._1554_ fd._1734_ fd._1719_ VGND VGND VPWR VPWR fd._1735_ sky130_fd_sc_hd__mux2_1
XFILLER_259_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5504_ fd._0375_ fd._0580_ VGND VGND VPWR VPWR fd._0581_ sky130_fd_sc_hd__xnor2_1
XFILLER_262_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6484_ fd._1648_ fd._1658_ VGND VGND VPWR VPWR fd._1659_ sky130_fd_sc_hd__nand2_1
XFILLER_140_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8223_ net71 net7 VGND VGND VPWR VPWR fd.a\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5435_ fd._0316_ VGND VGND VPWR VPWR fd._0506_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_283_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8154_ fd.a\[28\] fd.b\[28\] VGND VGND VPWR VPWR fd._3468_ sky130_fd_sc_hd__xnor2_1
XFILLER_55_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5366_ fd._0429_ VGND VGND VPWR VPWR fd._0430_ sky130_fd_sc_hd__clkinv_4
XFILLER_209_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_269_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7105_ fd._2340_ fd._2341_ VGND VGND VPWR VPWR fd._2343_ sky130_fd_sc_hd__xnor2_1
XFILLER_110_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4317_ fd._2573_ fd._2661_ fd._2639_ VGND VGND VPWR VPWR fd._2672_ sky130_fd_sc_hd__o21a_1
XFILLER_236_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8085_ fd._3409_ VGND VGND VPWR VPWR fd.mc\[10\] sky130_fd_sc_hd__clkbuf_1
Xfd._5297_ fd._0352_ fd._0353_ VGND VGND VPWR VPWR fd._0354_ sky130_fd_sc_hd__xor2_1
XFILLER_3_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7036_ fd._2076_ fd._2266_ VGND VGND VPWR VPWR fd._2267_ sky130_fd_sc_hd__and2_1
Xfd._4248_ fd._0362_ fd._0373_ VGND VGND VPWR VPWR fd._1913_ sky130_fd_sc_hd__xnor2_1
XFILLER_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4179_ fd._1143_ fd.a\[21\] VGND VGND VPWR VPWR fd._1154_ sky130_fd_sc_hd__and2_1
XFILLER_195_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_1675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7938_ fd._3258_ fd._3081_ VGND VGND VPWR VPWR fd._3259_ sky130_fd_sc_hd__nor2_1
XFILLER_164_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7869_ fd._2917_ fd._3182_ fd._3075_ VGND VGND VPWR VPWR fd._3183_ sky130_fd_sc_hd__mux2_1
XFILLER_117_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1468 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_276_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_269_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_265_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5220_ fd._0268_ VGND VGND VPWR VPWR fd._0269_ sky130_fd_sc_hd__buf_6
XTAP_5073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5151_ fd._4067_ fd._0067_ VGND VGND VPWR VPWR fd._0193_ sky130_fd_sc_hd__nand2_1
XTAP_4383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._4102_ fd._0296_ fd.a\[3\] VGND VGND VPWR VPWR fd._0307_ sky130_fd_sc_hd__or2_1
XTAP_3671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5082_ fd._4012_ fd._0116_ VGND VGND VPWR VPWR fd._0117_ sky130_fd_sc_hd__xnor2_1
XFILLER_75_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_257_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._5984_ fd._0541_ fd._1108_ VGND VGND VPWR VPWR fd._1109_ sky130_fd_sc_hd__nor2_1
XFILLER_146_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_277_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4935_ fd._3845_ VGND VGND VPWR VPWR fd._4029_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_185_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7723_ fd._2867_ fd._2851_ VGND VGND VPWR VPWR fd._3022_ sky130_fd_sc_hd__nor2_1
XFILLER_69_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7654_ fd._2377_ fd._2765_ VGND VGND VPWR VPWR fd._2946_ sky130_fd_sc_hd__nor2_1
Xfd._4866_ fd._3959_ VGND VGND VPWR VPWR fd._3960_ sky130_fd_sc_hd__buf_6
XFILLER_145_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_273_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6605_ fd._1789_ fd._1791_ fd._1720_ VGND VGND VPWR VPWR fd._1793_ sky130_fd_sc_hd__mux2_1
XFILLER_86_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_273_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7585_ fd._2665_ fd._2869_ VGND VGND VPWR VPWR fd._2871_ sky130_fd_sc_hd__or2_1
XFILLER_255_1668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4797_ fd._3667_ fd._3800_ VGND VGND VPWR VPWR fd._3891_ sky130_fd_sc_hd__nor2_1
XFILLER_259_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6536_ fd._1716_ VGND VGND VPWR VPWR fd._1717_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_87_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_259_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6467_ fd._1640_ fd._1622_ VGND VGND VPWR VPWR fd._1641_ sky130_fd_sc_hd__nor2_1
XFILLER_151_1644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5418_ fd._0486_ fd._0337_ VGND VGND VPWR VPWR fd._0487_ sky130_fd_sc_hd__xnor2_1
Xfd._8206_ net68 fd.ec\[7\] VGND VGND VPWR VPWR fd.c\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_151_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6398_ fd._1560_ fd._1564_ fd._1533_ VGND VGND VPWR VPWR fd._1565_ sky130_fd_sc_hd__mux2_1
XFILLER_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_283_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8137_ fd._3450_ fd._3451_ VGND VGND VPWR VPWR fd._3452_ sky130_fd_sc_hd__nor2_1
XFILLER_228_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5349_ fd._0409_ fd._0410_ VGND VGND VPWR VPWR fd._0411_ sky130_fd_sc_hd__nand2_1
XFILLER_215_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._8068_ fd._3077_ fd._3241_ fd._3398_ VGND VGND VPWR VPWR fd._3400_ sky130_fd_sc_hd__mux2_1
XFILLER_64_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7019_ fd._2032_ fd._2247_ fd._2021_ VGND VGND VPWR VPWR fd._2248_ sky130_fd_sc_hd__a21oi_1
XFILLER_35_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_260_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_278_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_278_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_262_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4720_ fd._3744_ fd._3741_ VGND VGND VPWR VPWR fd._3814_ sky130_fd_sc_hd__or2b_1
XFILLER_182_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_259_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4651_ fd._3738_ fd._3741_ fd._3743_ fd._3744_ VGND VGND VPWR VPWR fd._3745_ sky130_fd_sc_hd__a211o_1
XFILLER_155_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_1376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7370_ fd._2632_ fd._2633_ VGND VGND VPWR VPWR fd._2634_ sky130_fd_sc_hd__nor2_1
XFILLER_116_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4582_ fd._3535_ fd._3539_ VGND VGND VPWR VPWR fd._3676_ sky130_fd_sc_hd__or2_1
XFILLER_237_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_1688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_257_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6321_ fd._1278_ fd._1479_ fd._1422_ VGND VGND VPWR VPWR fd._1480_ sky130_fd_sc_hd__nand3b_1
XFILLER_2_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_256_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6252_ fd._1383_ fd._1390_ fd._1401_ fd._1402_ fd._1403_ VGND VGND VPWR VPWR fd._1404_
+ sky130_fd_sc_hd__a311o_1
XFILLER_2_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1606 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_266_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5203_ fd._0242_ fd._0244_ fd._0248_ fd._0249_ VGND VGND VPWR VPWR fd._0250_ sky130_fd_sc_hd__a211o_1
XFILLER_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6183_ fd._0768_ fd._1326_ VGND VGND VPWR VPWR fd._1328_ sky130_fd_sc_hd__and2_1
XFILLER_20_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_280_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5134_ fd._0172_ VGND VGND VPWR VPWR fd._0174_ sky130_fd_sc_hd__inv_2
XFILLER_209_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_252_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5065_ fd._3669_ fd._0096_ VGND VGND VPWR VPWR fd._0099_ sky130_fd_sc_hd__and2_1
XFILLER_221_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_15 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_222_1623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5967_ fd._0662_ fd._1086_ VGND VGND VPWR VPWR fd._1091_ sky130_fd_sc_hd__and2_1
XFILLER_161_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7706_ fd._3003_ VGND VGND VPWR VPWR fd._3004_ sky130_fd_sc_hd__clkinv_2
XFILLER_31_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_273_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4918_ fd._3689_ fd._3954_ fd._3958_ fd._4011_ VGND VGND VPWR VPWR fd._4012_ sky130_fd_sc_hd__a31o_1
XFILLER_133_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5898_ fd._0262_ VGND VGND VPWR VPWR fd._1015_ sky130_fd_sc_hd__buf_6
XFILLER_173_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_284_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4849_ fd._3035_ fd._3755_ fd._3757_ VGND VGND VPWR VPWR fd._3943_ sky130_fd_sc_hd__o21a_1
XFILLER_133_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7637_ fd._2141_ fd._2926_ VGND VGND VPWR VPWR fd._2928_ sky130_fd_sc_hd__nor2_1
XFILLER_115_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_255_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_170 VGND VGND VPWR VPWR user_project_wrapper_170/HI la_data_out[48]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_project_wrapper_181 VGND VGND VPWR VPWR user_project_wrapper_181/HI la_data_out[59]
+ sky130_fd_sc_hd__conb_1
Xuser_project_wrapper_192 VGND VGND VPWR VPWR user_project_wrapper_192/HI la_data_out[70]
+ sky130_fd_sc_hd__conb_1
XFILLER_82_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7568_ fd._2629_ fd._2659_ VGND VGND VPWR VPWR fd._2852_ sky130_fd_sc_hd__nand2_1
XFILLER_138_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6519_ fd._1494_ fd._1696_ VGND VGND VPWR VPWR fd._1698_ sky130_fd_sc_hd__nor2_1
XFILLER_134_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7499_ fd._2530_ fd._2775_ fd._2677_ VGND VGND VPWR VPWR fd._2776_ sky130_fd_sc_hd__mux2_1
XFILLER_5_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_284_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_284_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_270_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_221_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_9147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_267_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_247_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6870_ fd._1661_ fd._2013_ fd._2014_ VGND VGND VPWR VPWR fd._2084_ sky130_fd_sc_hd__mux2_1
XFILLER_141_1643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput13 io_in[20] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_2
XFILLER_278_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5821_ fd._0929_ VGND VGND VPWR VPWR fd._0930_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_200_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput24 io_in[30] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_1
XFILLER_15_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_1698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5752_ fd._0853_ fd._0777_ VGND VGND VPWR VPWR fd._0854_ sky130_fd_sc_hd__xnor2_1
XFILLER_115_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4703_ fd._3633_ fd._3749_ VGND VGND VPWR VPWR fd._3797_ sky130_fd_sc_hd__nand2_1
XFILLER_170_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5683_ fd._0771_ fd._0777_ VGND VGND VPWR VPWR fd._0778_ sky130_fd_sc_hd__nand2_1
XFILLER_131_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4634_ fd._3723_ fd.b\[12\] fd._3727_ VGND VGND VPWR VPWR fd._3728_ sky130_fd_sc_hd__mux2_1
Xfd._7422_ fd._2612_ fd._2690_ VGND VGND VPWR VPWR fd._2691_ sky130_fd_sc_hd__xnor2_1
XFILLER_112_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_285_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_258_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7353_ fd._1330_ fd._2508_ VGND VGND VPWR VPWR fd._2615_ sky130_fd_sc_hd__and2_1
XFILLER_123_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4565_ fd._3658_ fd._3502_ VGND VGND VPWR VPWR fd._3659_ sky130_fd_sc_hd__xnor2_1
XFILLER_285_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._6304_ fd._1263_ fd._1266_ VGND VGND VPWR VPWR fd._1461_ sky130_fd_sc_hd__or2_1
XFILLER_38_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7284_ fd._2380_ fd._2382_ VGND VGND VPWR VPWR fd._2539_ sky130_fd_sc_hd__and2_1
Xfd._4496_ fd._3588_ fd._3589_ VGND VGND VPWR VPWR fd._3590_ sky130_fd_sc_hd__nand2_1
XFILLER_211_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_244_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_285_1414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6235_ fd._0638_ fd._1210_ VGND VGND VPWR VPWR fd._1386_ sky130_fd_sc_hd__xnor2_1
XFILLER_96_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_253_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6166_ fd._1309_ fd._1078_ fd._1069_ VGND VGND VPWR VPWR fd._1310_ sky130_fd_sc_hd__o21bai_1
XFILLER_65_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5117_ fd._0091_ fd._0148_ fd._0154_ fd._0155_ VGND VGND VPWR VPWR fd._0156_ sky130_fd_sc_hd__a31o_1
XFILLER_209_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6097_ fd._1139_ fd._1138_ VGND VGND VPWR VPWR fd._1234_ sky130_fd_sc_hd__and2b_1
XFILLER_181_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_279_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5048_ fd._4019_ fd._4024_ fd._4026_ VGND VGND VPWR VPWR fd._0080_ sky130_fd_sc_hd__a21o_1
XFILLER_139_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6999_ fd._2225_ VGND VGND VPWR VPWR fd._2226_ sky130_fd_sc_hd__clkinv_4
XFILLER_146_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_276_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_264_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_275_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_8243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_8298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_273_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4350_ fd.b\[20\] VGND VGND VPWR VPWR fd._3035_ sky130_fd_sc_hd__buf_6
XFILLER_212_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_282_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_281_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4281_ fd.b\[9\] fd._2254_ VGND VGND VPWR VPWR fd._2276_ sky130_fd_sc_hd__nor2_1
XFILLER_47_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6020_ fd._0960_ fd._0964_ fd._0968_ VGND VGND VPWR VPWR fd._1149_ sky130_fd_sc_hd__o21ai_1
XFILLER_62_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_250_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7971_ fd._3152_ fd._3176_ VGND VGND VPWR VPWR fd._3295_ sky130_fd_sc_hd__nor2_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_28 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6922_ fd._1178_ VGND VGND VPWR VPWR fd._2141_ sky130_fd_sc_hd__buf_6
XFILLER_147_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6853_ fd._1856_ fd._2064_ fd._2020_ VGND VGND VPWR VPWR fd._2065_ sky130_fd_sc_hd__mux2_1
XFILLER_163_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5804_ fd._0676_ fd._0688_ VGND VGND VPWR VPWR fd._0911_ sky130_fd_sc_hd__nand2_1
XFILLER_129_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6784_ fd._1743_ fd._1988_ fd._1917_ VGND VGND VPWR VPWR fd._1989_ sky130_fd_sc_hd__mux2_1
XFILLER_116_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5735_ fd._0826_ fd._0831_ fd._0833_ fd._0834_ VGND VGND VPWR VPWR fd._0836_ sky130_fd_sc_hd__a31o_1
XFILLER_171_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5666_ fd._0592_ fd._0759_ VGND VGND VPWR VPWR fd._0760_ sky130_fd_sc_hd__nand2_1
XFILLER_217_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4617_ fd._0857_ fd._3650_ VGND VGND VPWR VPWR fd._3711_ sky130_fd_sc_hd__and2_1
Xfd._7405_ fd._2503_ fd._2671_ fd._2472_ VGND VGND VPWR VPWR fd._2673_ sky130_fd_sc_hd__o21ai_1
XFILLER_217_1588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5597_ fd._0644_ VGND VGND VPWR VPWR fd._0684_ sky130_fd_sc_hd__inv_2
XFILLER_150_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4548_ fd.b\[14\] fd._3310_ fd._3449_ fd._3641_ VGND VGND VPWR VPWR fd._3642_
+ sky130_fd_sc_hd__o2bb2a_1
Xfd._7336_ fd._2399_ fd._2403_ VGND VGND VPWR VPWR fd._2597_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7267_ fd._2519_ fd._2520_ VGND VGND VPWR VPWR fd._2521_ sky130_fd_sc_hd__xor2_1
XFILLER_285_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._4479_ fd._3572_ VGND VGND VPWR VPWR fd._3573_ sky130_fd_sc_hd__inv_2
XFILLER_214_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_285_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6218_ fd._1364_ fd._1366_ VGND VGND VPWR VPWR fd._1367_ sky130_fd_sc_hd__xnor2_1
XFILLER_26_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_246_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7198_ fd._1330_ fd._2443_ VGND VGND VPWR VPWR fd._2445_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_253_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6149_ fd._1290_ fd._1237_ VGND VGND VPWR VPWR fd._1291_ sky130_fd_sc_hd__and2_1
XFILLER_213_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_257_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_1579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_1570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_1579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_263_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_264_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_8051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5520_ fd._0282_ fd._0598_ VGND VGND VPWR VPWR fd._0599_ sky130_fd_sc_hd__xnor2_1
XFILLER_193_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5451_ fd._0427_ fd._0426_ VGND VGND VPWR VPWR fd._0523_ sky130_fd_sc_hd__nor2_1
XFILLER_136_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4402_ fd._2155_ fd._3495_ VGND VGND VPWR VPWR fd._3496_ sky130_fd_sc_hd__or2_1
XTAP_6671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._8170_ fd._3483_ fd._3484_ VGND VGND VPWR VPWR fd.ec\[6\] sky130_fd_sc_hd__nand2_1
XFILLER_136_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._5382_ fd._0436_ fd._0443_ fd._0445_ fd._0446_ VGND VGND VPWR VPWR fd._0447_ sky130_fd_sc_hd__a31o_1
XTAP_6693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_255_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_282_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7121_ fd._1559_ fd._2359_ VGND VGND VPWR VPWR fd._2360_ sky130_fd_sc_hd__nand2_1
Xfd._4333_ fd._0109_ fd._2837_ fd._0032_ VGND VGND VPWR VPWR fd._2848_ sky130_fd_sc_hd__o21bai_1
XFILLER_181_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7052_ fd._2278_ fd._2283_ VGND VGND VPWR VPWR fd._2284_ sky130_fd_sc_hd__nor2_1
XFILLER_63_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4264_ fd._1660_ fd._0241_ fd._0263_ fd._0472_ VGND VGND VPWR VPWR fd._2089_ sky130_fd_sc_hd__o31a_1
XFILLER_169_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6003_ fd._0953_ fd._1129_ fd._1046_ VGND VGND VPWR VPWR fd._1130_ sky130_fd_sc_hd__and3_1
XFILLER_169_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4195_ fd._1319_ VGND VGND VPWR VPWR fd._1330_ sky130_fd_sc_hd__buf_6
XFILLER_23_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7954_ fd._2763_ fd._3265_ fd._3274_ VGND VGND VPWR VPWR fd._3276_ sky130_fd_sc_hd__o21a_1
XFILLER_108_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6905_ fd._2119_ fd._2120_ fd._2116_ fd._2121_ VGND VGND VPWR VPWR fd._2123_ sky130_fd_sc_hd__a31o_1
XFILLER_148_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_1592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7885_ fd._3110_ fd._3111_ VGND VGND VPWR VPWR fd._3201_ sky130_fd_sc_hd__nor2_1
XFILLER_163_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6836_ fd._2021_ fd._2046_ VGND VGND VPWR VPWR fd._2047_ sky130_fd_sc_hd__nand2_1
XFILLER_239_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6767_ fd._1970_ fd._1813_ VGND VGND VPWR VPWR fd._1971_ sky130_fd_sc_hd__nand2_1
XFILLER_171_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5718_ fd._0427_ fd._0816_ VGND VGND VPWR VPWR fd._0817_ sky130_fd_sc_hd__nor2_1
XFILLER_67_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6698_ fd._1319_ fd._1894_ VGND VGND VPWR VPWR fd._1895_ sky130_fd_sc_hd__nor2_1
XFILLER_277_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._5649_ fd._0572_ fd._0740_ VGND VGND VPWR VPWR fd._0741_ sky130_fd_sc_hd__xor2_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7319_ fd._2396_ fd._2568_ fd._2345_ VGND VGND VPWR VPWR fd._2578_ sky130_fd_sc_hd__a21boi_1
XFILLER_79_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_253_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_1492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_268_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_277_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_242_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4951_ fd._3914_ fd._4044_ fd._3960_ VGND VGND VPWR VPWR fd._4045_ sky130_fd_sc_hd__mux2_1
XFILLER_125_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4882_ fd._3708_ fd._3892_ VGND VGND VPWR VPWR fd._3976_ sky130_fd_sc_hd__and2_1
Xfd._7670_ fd._0312_ fd._2935_ fd._2944_ fd._2962_ fd._2963_ VGND VGND VPWR VPWR fd._2964_
+ sky130_fd_sc_hd__a221o_1
XFILLER_177_1620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_246_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6621_ fd._1618_ fd._1809_ VGND VGND VPWR VPWR fd._1810_ sky130_fd_sc_hd__nand2_1
XFILLER_177_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6552_ fd._1557_ fd._1733_ VGND VGND VPWR VPWR fd._1734_ sky130_fd_sc_hd__xnor2_1
XFILLER_158_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_259_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_1552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5503_ fd._0385_ fd._0379_ VGND VGND VPWR VPWR fd._0580_ sky130_fd_sc_hd__and2b_1
Xfd._6483_ fd._1650_ fd._1655_ fd._1657_ VGND VGND VPWR VPWR fd._1658_ sky130_fd_sc_hd__a21oi_1
XFILLER_45_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8222_ net71 net6 VGND VGND VPWR VPWR fd.a\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_136_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5434_ fd._3669_ VGND VGND VPWR VPWR fd._0504_ sky130_fd_sc_hd__buf_6
XFILLER_214_1558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_267_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_283_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5365_ fd._0427_ fd._0426_ VGND VGND VPWR VPWR fd._0429_ sky130_fd_sc_hd__xnor2_1
Xfd._8153_ fd._3466_ fd._3467_ VGND VGND VPWR VPWR fd.ec\[4\] sky130_fd_sc_hd__nand2_1
XFILLER_94_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4316_ fd._2639_ fd._2650_ VGND VGND VPWR VPWR fd._2661_ sky130_fd_sc_hd__nand2_1
Xfd._7104_ fd._2140_ fd._2193_ VGND VGND VPWR VPWR fd._2341_ sky130_fd_sc_hd__and2b_1
XFILLER_48_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5296_ fd._0155_ fd._0154_ VGND VGND VPWR VPWR fd._0353_ sky130_fd_sc_hd__or2b_1
Xfd._8084_ fd._1617_ fd._1813_ fd._3398_ VGND VGND VPWR VPWR fd._3409_ sky130_fd_sc_hd__mux2_1
XFILLER_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_282_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_235_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4247_ fd.a\[1\] VGND VGND VPWR VPWR fd._1902_ sky130_fd_sc_hd__clkinv_2
Xfd._7035_ fd._2087_ fd._2264_ fd._2116_ VGND VGND VPWR VPWR fd._2266_ sky130_fd_sc_hd__mux2_1
XFILLER_251_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._4178_ fd.b\[21\] VGND VGND VPWR VPWR fd._1143_ sky130_fd_sc_hd__inv_2
XFILLER_251_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_1643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7937_ fd._3080_ VGND VGND VPWR VPWR fd._3258_ sky130_fd_sc_hd__inv_2
XFILLER_109_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7868_ fd._2975_ fd._3181_ VGND VGND VPWR VPWR fd._3182_ sky130_fd_sc_hd__xor2_1
XTAP_8809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6819_ fd._2027_ fd._1832_ fd._1820_ VGND VGND VPWR VPWR fd._2028_ sky130_fd_sc_hd__a21o_1
XFILLER_102_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7799_ fd._2977_ fd._2984_ fd._2987_ VGND VGND VPWR VPWR fd._3106_ sky130_fd_sc_hd__a21o_1
XFILLER_258_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_1606 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_277_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_252_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_285_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_226_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_277_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_265_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_264_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5150_ fd._4069_ fd._4068_ fd._4062_ VGND VGND VPWR VPWR fd._0192_ sky130_fd_sc_hd__a21oi_1
XTAP_4373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4101_ fd.b\[3\] VGND VGND VPWR VPWR fd._0296_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_218_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5081_ fd._0115_ fd._4010_ VGND VGND VPWR VPWR fd._0116_ sky130_fd_sc_hd__or2_1
XFILLER_233_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5983_ fd._0938_ fd._1107_ fd._1046_ VGND VGND VPWR VPWR fd._1108_ sky130_fd_sc_hd__mux2_1
XFILLER_257_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7722_ fd._2465_ fd._3019_ fd._3020_ VGND VGND VPWR VPWR fd._3021_ sky130_fd_sc_hd__mux2_1
XFILLER_9_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4934_ fd._4019_ fd._4024_ fd._4025_ fd._4026_ fd._4027_ VGND VGND VPWR VPWR fd._4028_
+ sky130_fd_sc_hd__a2111o_1
XFILLER_145_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_255_1603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._7653_ fd._2759_ fd._2762_ VGND VGND VPWR VPWR fd._2945_ sky130_fd_sc_hd__or2_1
Xfd._4865_ fd._3954_ fd._3958_ VGND VGND VPWR VPWR fd._3959_ sky130_fd_sc_hd__nand2_4
XFILLER_161_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_255_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._6604_ fd._1790_ fd._1606_ VGND VGND VPWR VPWR fd._1791_ sky130_fd_sc_hd__xor2_1
Xfd._7584_ fd._2863_ fd._2667_ fd._2853_ VGND VGND VPWR VPWR fd._2869_ sky130_fd_sc_hd__o21a_1
XFILLER_113_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4796_ fd._3674_ fd._3701_ fd._3671_ VGND VGND VPWR VPWR fd._3890_ sky130_fd_sc_hd__o21ai_1
XFILLER_114_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6535_ fd._0131_ fd._1714_ VGND VGND VPWR VPWR fd._1716_ sky130_fd_sc_hd__nor2_1
XFILLER_64_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_256_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_253_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6466_ fd._2738_ fd._1639_ VGND VGND VPWR VPWR fd._1640_ sky130_fd_sc_hd__nor2_1
XFILLER_25_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8205_ net68 fd.ec\[6\] VGND VGND VPWR VPWR fd.c\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_267_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5417_ fd._0341_ fd._0485_ fd._0301_ VGND VGND VPWR VPWR fd._0486_ sky130_fd_sc_hd__o21ai_1
XFILLER_283_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6397_ fd._1562_ fd._1563_ VGND VGND VPWR VPWR fd._1564_ sky130_fd_sc_hd__xnor2_1
XFILLER_56_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8136_ fd.a\[26\] fd.b\[26\] VGND VGND VPWR VPWR fd._3451_ sky130_fd_sc_hd__and2b_1
XFILLER_283_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5348_ fd._0026_ fd._0408_ VGND VGND VPWR VPWR fd._0410_ sky130_fd_sc_hd__nand2_1
XFILLER_3_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5279_ fd._0096_ fd._0269_ VGND VGND VPWR VPWR fd._0334_ sky130_fd_sc_hd__nor2_1
XFILLER_222_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8067_ fd._3399_ VGND VGND VPWR VPWR fd.mc\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_24_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7018_ fd._2246_ fd._2046_ fd._2026_ VGND VGND VPWR VPWR fd._2247_ sky130_fd_sc_hd__a21o_1
XFILLER_145_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_223_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_225_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_28 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_258_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_1583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_278_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_259_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_263_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_262_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_265_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_262_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_259_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4650_ fd._1297_ fd._3740_ VGND VGND VPWR VPWR fd._3744_ sky130_fd_sc_hd__and2_1
XFILLER_100_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._4581_ fd._0219_ VGND VGND VPWR VPWR fd._3675_ sky130_fd_sc_hd__buf_6
XFILLER_9_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6320_ fd._1118_ fd._1277_ VGND VGND VPWR VPWR fd._1479_ sky130_fd_sc_hd__nand2_1
XFILLER_123_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6251_ fd._0807_ fd._1376_ VGND VGND VPWR VPWR fd._1403_ sky130_fd_sc_hd__nor2_1
XFILLER_250_1588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5202_ fd._0126_ fd._0245_ fd._0247_ VGND VGND VPWR VPWR fd._0249_ sky130_fd_sc_hd__a21oi_1
XFILLER_225_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6182_ fd._0768_ fd._1326_ VGND VGND VPWR VPWR fd._1327_ sky130_fd_sc_hd__nor2_1
XFILLER_266_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_264_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5133_ fd._3917_ fd._0172_ VGND VGND VPWR VPWR fd._0173_ sky130_fd_sc_hd__or2_1
XFILLER_111_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_252_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_280_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5064_ fd._3669_ fd._0096_ VGND VGND VPWR VPWR fd._0097_ sky130_fd_sc_hd__nor2_1
XFILLER_127_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_16 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_277_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5966_ fd._1083_ fd._1087_ fd._1089_ VGND VGND VPWR VPWR fd._1090_ sky130_fd_sc_hd__o21a_1
XFILLER_146_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._7705_ fd._2999_ fd._3001_ VGND VGND VPWR VPWR fd._3003_ sky130_fd_sc_hd__xnor2_1
Xfd._4917_ fd.b\[1\] VGND VGND VPWR VPWR fd._4011_ sky130_fd_sc_hd__buf_6
XFILLER_146_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5897_ fd._0450_ fd._1013_ VGND VGND VPWR VPWR fd._1014_ sky130_fd_sc_hd__xnor2_2
XFILLER_12_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7636_ fd._2141_ fd._2926_ VGND VGND VPWR VPWR fd._2927_ sky130_fd_sc_hd__and2_1
Xfd._4848_ fd._3795_ fd._3935_ fd._3939_ VGND VGND VPWR VPWR fd._3942_ sky130_fd_sc_hd__a21o_1
XFILLER_161_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_project_wrapper_160 VGND VGND VPWR VPWR user_project_wrapper_160/HI la_data_out[38]
+ sky130_fd_sc_hd__conb_1
XFILLER_82_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_171 VGND VGND VPWR VPWR user_project_wrapper_171/HI la_data_out[49]
+ sky130_fd_sc_hd__conb_1
XFILLER_88_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_project_wrapper_182 VGND VGND VPWR VPWR user_project_wrapper_182/HI la_data_out[60]
+ sky130_fd_sc_hd__conb_1
XFILLER_86_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_255_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7567_ fd._2816_ fd._2819_ fd._2830_ fd._2847_ fd._2850_ VGND VGND VPWR VPWR fd._2851_
+ sky130_fd_sc_hd__o311a_1
Xuser_project_wrapper_193 VGND VGND VPWR VPWR user_project_wrapper_193/HI la_data_out[71]
+ sky130_fd_sc_hd__conb_1
XFILLER_276_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4779_ fd._3872_ fd._3693_ fd._3786_ VGND VGND VPWR VPWR fd._3873_ sky130_fd_sc_hd__mux2_1
XFILLER_141_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6518_ fd._1494_ fd._1696_ VGND VGND VPWR VPWR fd._1697_ sky130_fd_sc_hd__nand2_1
XFILLER_29_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7498_ fd._2531_ fd._2774_ VGND VGND VPWR VPWR fd._2775_ sky130_fd_sc_hd__xnor2_1
XFILLER_64_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6449_ fd._1510_ fd._1620_ fd._1615_ VGND VGND VPWR VPWR fd._1621_ sky130_fd_sc_hd__mux2_1
XFILLER_56_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8119_ fd._3432_ fd._3433_ VGND VGND VPWR VPWR fd._3434_ sky130_fd_sc_hd__nor2_1
XFILLER_270_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_1551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_270_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1634 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_9148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_273_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_1675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1635 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput14 io_in[21] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_4
XFILLER_204_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5820_ fd._0928_ fd._0922_ VGND VGND VPWR VPWR fd._0929_ sky130_fd_sc_hd__nor2_1
XFILLER_174_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput25 io_in[31] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_1
XFILLER_278_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5751_ fd._0851_ fd._0852_ fd._0767_ VGND VGND VPWR VPWR fd._0853_ sky130_fd_sc_hd__o21ai_1
XFILLER_183_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4702_ fd._3637_ fd._3748_ VGND VGND VPWR VPWR fd._3796_ sky130_fd_sc_hd__nand2_1
Xfd._5682_ fd._0775_ fd._0776_ VGND VGND VPWR VPWR fd._0777_ sky130_fd_sc_hd__and2_1
XFILLER_170_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_254_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7421_ fd._2677_ fd._2689_ VGND VGND VPWR VPWR fd._2690_ sky130_fd_sc_hd__nand2_1
Xfd._4633_ fd._1451_ fd._3726_ VGND VGND VPWR VPWR fd._3727_ sky130_fd_sc_hd__xnor2_1
XFILLER_130_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_252_1639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._7352_ fd._2076_ fd._2608_ fd._2613_ VGND VGND VPWR VPWR fd._2614_ sky130_fd_sc_hd__mux2_1
Xfd._4564_ fd._0428_ VGND VGND VPWR VPWR fd._3658_ sky130_fd_sc_hd__clkinv_2
XFILLER_170_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_257_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6303_ fd._1255_ VGND VGND VPWR VPWR fd._1460_ sky130_fd_sc_hd__clkinv_2
XFILLER_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_285_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_266_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4495_ fd.b\[19\] fd._3587_ VGND VGND VPWR VPWR fd._3589_ sky130_fd_sc_hd__or2_1
XFILLER_211_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7283_ fd._2533_ fd._2537_ VGND VGND VPWR VPWR fd._2538_ sky130_fd_sc_hd__nand2_1
XFILLER_38_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_272_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6234_ fd._1211_ fd._1206_ VGND VGND VPWR VPWR fd._1384_ sky130_fd_sc_hd__nand2_1
XFILLER_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6165_ fd._1162_ fd._1166_ VGND VGND VPWR VPWR fd._1309_ sky130_fd_sc_hd__nand2_1
XFILLER_20_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_279_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5116_ fd._3905_ fd._0152_ VGND VGND VPWR VPWR fd._0155_ sky130_fd_sc_hd__and2_1
Xfd._6096_ fd._1229_ fd._1230_ fd._1232_ VGND VGND VPWR VPWR fd._1233_ sky130_fd_sc_hd__mux2_1
XFILLER_20_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5047_ fd._0078_ fd._4040_ fd._0060_ VGND VGND VPWR VPWR fd._0079_ sky130_fd_sc_hd__mux2_1
XFILLER_221_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6998_ fd._2223_ fd._2224_ VGND VGND VPWR VPWR fd._2225_ sky130_fd_sc_hd__and2_1
XFILLER_147_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5949_ fd._1070_ fd._1052_ VGND VGND VPWR VPWR fd._1071_ sky130_fd_sc_hd__nand2_1
XFILLER_107_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7619_ fd._2906_ fd._2907_ VGND VGND VPWR VPWR fd._2908_ sky130_fd_sc_hd__nor2_1
XTAP_6319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_276_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1550 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_276_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_249_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_249_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_1376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_1576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_275_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_8222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_8233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_279_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_251_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_281_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4280_ fd.b\[9\] fd._2254_ VGND VGND VPWR VPWR fd._2265_ sky130_fd_sc_hd__nand2_1
XFILLER_267_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_267_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_263_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7970_ fd._2142_ fd._3158_ fd._3175_ VGND VGND VPWR VPWR fd._3294_ sky130_fd_sc_hd__a21o_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6921_ fd._2135_ fd._2139_ VGND VGND VPWR VPWR fd._2140_ sky130_fd_sc_hd__nor2_1
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6852_ fd._1685_ fd._1898_ VGND VGND VPWR VPWR fd._2064_ sky130_fd_sc_hd__xnor2_1
XFILLER_15_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5803_ fd._0909_ VGND VGND VPWR VPWR fd._0910_ sky130_fd_sc_hd__inv_2
XFILLER_200_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6783_ fd._1926_ fd._1987_ VGND VGND VPWR VPWR fd._1988_ sky130_fd_sc_hd__nor2_1
XFILLER_265_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5734_ fd._0262_ fd._0825_ VGND VGND VPWR VPWR fd._0834_ sky130_fd_sc_hd__nor2_1
XFILLER_274_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5665_ fd._0594_ fd._0757_ VGND VGND VPWR VPWR fd._0759_ sky130_fd_sc_hd__xnor2_1
XFILLER_135_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7404_ fd._2662_ fd._2479_ fd._2477_ VGND VGND VPWR VPWR fd._2671_ sky130_fd_sc_hd__a21oi_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4616_ fd._3702_ fd._3705_ fd._3707_ fd._3709_ VGND VGND VPWR VPWR fd._3710_ sky130_fd_sc_hd__a211o_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5596_ fd._0682_ VGND VGND VPWR VPWR fd._0683_ sky130_fd_sc_hd__inv_2
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_258_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7335_ fd._2586_ fd._2594_ fd._2591_ VGND VGND VPWR VPWR fd._2596_ sky130_fd_sc_hd__o21ai_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4547_ fd._3439_ fd._3640_ fd._3376_ VGND VGND VPWR VPWR fd._3641_ sky130_fd_sc_hd__o21ai_1
XFILLER_135_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_257_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_285_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._7266_ fd._2360_ fd._2387_ VGND VGND VPWR VPWR fd._2520_ sky130_fd_sc_hd__nand2_1
XFILLER_113_1554 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4478_ fd.b\[17\] fd._3571_ VGND VGND VPWR VPWR fd._3572_ sky130_fd_sc_hd__xnor2_1
XFILLER_211_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6217_ fd._1189_ fd._1365_ VGND VGND VPWR VPWR fd._1366_ sky130_fd_sc_hd__nand2_1
XFILLER_93_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7197_ fd._1330_ fd._2443_ VGND VGND VPWR VPWR fd._2444_ sky130_fd_sc_hd__or2_1
XFILLER_81_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_281_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6148_ fd._0965_ fd._1236_ VGND VGND VPWR VPWR fd._1290_ sky130_fd_sc_hd__nand2_1
XFILLER_230_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_1516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6079_ fd._0450_ fd._1195_ VGND VGND VPWR VPWR fd._1214_ sky130_fd_sc_hd__and2_1
XFILLER_34_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_263_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_270_1558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_1678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_260_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_1627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_279_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5450_ fd._3883_ fd._0518_ VGND VGND VPWR VPWR fd._0522_ sky130_fd_sc_hd__nor2_1
XFILLER_80_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4401_ fd._2111_ fd._3494_ fd._3211_ VGND VGND VPWR VPWR fd._3495_ sky130_fd_sc_hd__mux2_1
XFILLER_132_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5381_ fd._0262_ fd._0435_ VGND VGND VPWR VPWR fd._0446_ sky130_fd_sc_hd__nor2_1
XTAP_6683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7120_ fd._2356_ fd._2358_ fd._2322_ VGND VGND VPWR VPWR fd._2359_ sky130_fd_sc_hd__mux2_1
XFILLER_282_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4332_ fd._0054_ fd._2826_ VGND VGND VPWR VPWR fd._2837_ sky130_fd_sc_hd__nor2_1
XTAP_5982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7051_ fd._2098_ fd._2282_ fd._2116_ VGND VGND VPWR VPWR fd._2283_ sky130_fd_sc_hd__mux2_1
Xfd._4263_ fd._1759_ fd._2056_ fd._2067_ VGND VGND VPWR VPWR fd._2078_ sky130_fd_sc_hd__a21oi_1
XFILLER_47_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6002_ fd._1118_ fd._0903_ fd._0952_ VGND VGND VPWR VPWR fd._1129_ sky130_fd_sc_hd__nand3_1
XFILLER_282_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4194_ fd._1308_ VGND VGND VPWR VPWR fd._1319_ sky130_fd_sc_hd__buf_6
XFILLER_63_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7953_ fd._2763_ fd._1970_ VGND VGND VPWR VPWR fd._3275_ sky130_fd_sc_hd__or2_1
XFILLER_128_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6904_ fd._2009_ fd._2116_ VGND VGND VPWR VPWR fd._2121_ sky130_fd_sc_hd__nor2_1
XFILLER_108_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7884_ fd._3116_ fd._3198_ VGND VGND VPWR VPWR fd._3199_ sky130_fd_sc_hd__nor2_1
XFILLER_258_1612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6835_ fd._2738_ fd._2025_ VGND VGND VPWR VPWR fd._2046_ sky130_fd_sc_hd__xnor2_1
XFILLER_159_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_258_1634 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_278_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6766_ fd._0437_ VGND VGND VPWR VPWR fd._1970_ sky130_fd_sc_hd__buf_6
XFILLER_116_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5717_ fd._0629_ fd._0815_ fd._0801_ VGND VGND VPWR VPWR fd._0816_ sky130_fd_sc_hd__mux2_1
XFILLER_171_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6697_ fd._1672_ fd._1893_ fd._1720_ VGND VGND VPWR VPWR fd._1894_ sky130_fd_sc_hd__mux2_1
XFILLER_132_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5648_ fd._0578_ fd._0577_ VGND VGND VPWR VPWR fd._0740_ sky130_fd_sc_hd__and2b_1
XFILLER_63_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5579_ fd._0525_ fd._0663_ VGND VGND VPWR VPWR fd._0664_ sky130_fd_sc_hd__xnor2_1
XFILLER_273_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7318_ fd._2506_ VGND VGND VPWR VPWR fd._2577_ sky130_fd_sc_hd__inv_6
XFILLER_6_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7249_ fd._2469_ fd._2316_ fd._2245_ VGND VGND VPWR VPWR fd._2501_ sky130_fd_sc_hd__a21o_1
XFILLER_26_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_263_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_269_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_1495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_246_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4950_ fd._3908_ fd._4043_ VGND VGND VPWR VPWR fd._4044_ sky130_fd_sc_hd__xnor2_1
XFILLER_199_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4881_ fd._3850_ fd._3974_ fd._3959_ VGND VGND VPWR VPWR fd._3975_ sky130_fd_sc_hd__mux2_1
XFILLER_8_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6620_ fd._1622_ fd._1808_ VGND VGND VPWR VPWR fd._1809_ sky130_fd_sc_hd__or2_1
XFILLER_275_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6551_ fd._1566_ fd._1596_ VGND VGND VPWR VPWR fd._1733_ sky130_fd_sc_hd__and2_1
XFILLER_153_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_271_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5502_ fd._0572_ fd._0577_ fd._0578_ VGND VGND VPWR VPWR fd._0579_ sky130_fd_sc_hd__a21oi_1
XFILLER_49_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._6482_ fd._1656_ fd._1654_ VGND VGND VPWR VPWR fd._1657_ sky130_fd_sc_hd__nor2_1
XFILLER_262_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8221_ net71 net5 VGND VGND VPWR VPWR fd.a\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_7192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5433_ fd._0496_ fd._0501_ fd._0502_ VGND VGND VPWR VPWR fd._0503_ sky130_fd_sc_hd__a21o_1
XFILLER_136_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8152_ fd._3456_ fd._3465_ VGND VGND VPWR VPWR fd._3467_ sky130_fd_sc_hd__or2_1
Xfd._5364_ fd._3675_ VGND VGND VPWR VPWR fd._0427_ sky130_fd_sc_hd__buf_6
XFILLER_132_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_282_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7103_ fd._2151_ fd._2158_ fd._2192_ fd._2194_ VGND VGND VPWR VPWR fd._2340_ sky130_fd_sc_hd__o31a_1
XFILLER_3_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4315_ fd._2584_ fd._2628_ VGND VGND VPWR VPWR fd._2650_ sky130_fd_sc_hd__nand2_1
XFILLER_283_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8083_ fd._3408_ VGND VGND VPWR VPWR fd.mc\[9\] sky130_fd_sc_hd__clkbuf_1
XFILLER_282_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5295_ fd._0091_ fd._0148_ VGND VGND VPWR VPWR fd._0352_ sky130_fd_sc_hd__nand2_1
XFILLER_48_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7034_ fd._2084_ fd._2263_ VGND VGND VPWR VPWR fd._2264_ sky130_fd_sc_hd__xnor2_1
Xfd._4246_ fd.b\[3\] fd._1880_ VGND VGND VPWR VPWR fd._1891_ sky130_fd_sc_hd__nand2_1
XFILLER_235_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4177_ fd._0175_ fd._1077_ fd._1121_ VGND VGND VPWR VPWR fd._1132_ sky130_fd_sc_hd__a21oi_1
XFILLER_225_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_251_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7936_ fd._3087_ fd._3212_ VGND VGND VPWR VPWR fd._3257_ sky130_fd_sc_hd__or2_1
XFILLER_17_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7867_ fd._2965_ fd._2971_ fd._2973_ VGND VGND VPWR VPWR fd._3181_ sky130_fd_sc_hd__a21oi_1
XFILLER_164_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6818_ fd._2018_ VGND VGND VPWR VPWR fd._2027_ sky130_fd_sc_hd__inv_2
XFILLER_117_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7798_ fd._3099_ fd._3103_ fd._3104_ VGND VGND VPWR VPWR fd._3105_ sky130_fd_sc_hd__a21o_1
XFILLER_258_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6749_ fd._1767_ fd._1772_ VGND VGND VPWR VPWR fd._1951_ sky130_fd_sc_hd__nand2_1
XFILLER_172_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_252_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_259_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_274_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_277_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_264_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4100_ fd._0230_ fd._0274_ VGND VGND VPWR VPWR fd._0285_ sky130_fd_sc_hd__nand2_1
XTAP_4396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5080_ fd._3688_ fd._0114_ VGND VGND VPWR VPWR fd._0115_ sky130_fd_sc_hd__nor2_1
XFILLER_40_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_281_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5982_ fd._1105_ fd._1106_ VGND VGND VPWR VPWR fd._1107_ sky130_fd_sc_hd__xnor2_1
XFILLER_125_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7721_ fd._0131_ fd._2879_ VGND VGND VPWR VPWR fd._3020_ sky130_fd_sc_hd__xnor2_2
Xfd._4933_ fd._2155_ fd._3979_ VGND VGND VPWR VPWR fd._4027_ sky130_fd_sc_hd__xnor2_1
XFILLER_220_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7652_ fd._2942_ fd._2943_ VGND VGND VPWR VPWR fd._2944_ sky130_fd_sc_hd__and2_1
Xfd._4864_ fd._3947_ fd._3946_ fd._3949_ fd._3957_ VGND VGND VPWR VPWR fd._3958_ sky130_fd_sc_hd__o31a_2
XFILLER_138_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6603_ fd._1543_ fd._1779_ fd._1541_ VGND VGND VPWR VPWR fd._1790_ sky130_fd_sc_hd__a21bo_1
XFILLER_275_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7583_ fd._2867_ fd._2866_ VGND VGND VPWR VPWR fd._2868_ sky130_fd_sc_hd__and2_1
Xfd._4795_ fd._3671_ fd._3674_ fd._3701_ VGND VGND VPWR VPWR fd._3889_ sky130_fd_sc_hd__or3_1
XFILLER_259_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6534_ fd._1708_ VGND VGND VPWR VPWR fd._1714_ sky130_fd_sc_hd__inv_2
XFILLER_138_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_259_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6465_ fd._1621_ VGND VGND VPWR VPWR fd._1639_ sky130_fd_sc_hd__inv_2
XFILLER_101_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8204_ net68 fd.ec\[5\] VGND VGND VPWR VPWR fd.c\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_25_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5416_ fd._0330_ fd._0336_ fd._0338_ VGND VGND VPWR VPWR fd._0485_ sky130_fd_sc_hd__a21o_1
XFILLER_56_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_267_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6396_ fd._1390_ fd._1401_ VGND VGND VPWR VPWR fd._1563_ sky130_fd_sc_hd__nand2_1
XFILLER_3_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_249_1408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8135_ fd.b\[26\] fd.a\[26\] VGND VGND VPWR VPWR fd._3450_ sky130_fd_sc_hd__and2b_1
XFILLER_186_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._5347_ fd._0026_ fd._0408_ VGND VGND VPWR VPWR fd._0409_ sky130_fd_sc_hd__or2_1
XFILLER_243_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1580 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8066_ fd._3241_ fd._3395_ fd._3398_ VGND VGND VPWR VPWR fd._3399_ sky130_fd_sc_hd__mux2_4
XFILLER_64_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5278_ fd._0100_ fd._0331_ VGND VGND VPWR VPWR fd._0333_ sky130_fd_sc_hd__or2_1
XFILLER_110_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7017_ fd._2236_ VGND VGND VPWR VPWR fd._2246_ sky130_fd_sc_hd__inv_2
Xfd._4229_ fd.b\[6\] fd._1693_ VGND VGND VPWR VPWR fd._1704_ sky130_fd_sc_hd__and2_1
XFILLER_251_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_260_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7919_ fd._3026_ fd._3237_ VGND VGND VPWR VPWR fd._3238_ sky130_fd_sc_hd__xnor2_1
XFILLER_109_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_258_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_278_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_1558 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_272_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_269_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4580_ fd._0252_ fd._3673_ VGND VGND VPWR VPWR fd._3674_ sky130_fd_sc_hd__and2_1
XFILLER_155_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_257_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_1523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6250_ fd._0450_ fd._1382_ VGND VGND VPWR VPWR fd._1402_ sky130_fd_sc_hd__and2_1
XFILLER_133_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5201_ fd._0126_ fd._0245_ fd._0247_ VGND VGND VPWR VPWR fd._0248_ sky130_fd_sc_hd__and3_1
XFILLER_77_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6181_ fd._1164_ fd._1325_ VGND VGND VPWR VPWR fd._1326_ sky130_fd_sc_hd__xnor2_1
XFILLER_168_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1690 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5132_ fd._4045_ fd._0061_ fd._0171_ VGND VGND VPWR VPWR fd._0172_ sky130_fd_sc_hd__o21ai_1
XTAP_4193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._5063_ fd._0095_ fd._3992_ fd._0059_ VGND VGND VPWR VPWR fd._0096_ sky130_fd_sc_hd__mux2_1
XFILLER_233_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_17 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5965_ fd._0916_ fd._1082_ VGND VGND VPWR VPWR fd._1089_ sky130_fd_sc_hd__nand2_1
XFILLER_186_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4916_ fd._4006_ fd._4009_ fd._3688_ VGND VGND VPWR VPWR fd._4010_ sky130_fd_sc_hd__o21a_1
XFILLER_179_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._7704_ fd._3000_ fd._2802_ VGND VGND VPWR VPWR fd._3001_ sky130_fd_sc_hd__nor2_1
XFILLER_277_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5896_ fd._0825_ fd._1012_ fd._0998_ VGND VGND VPWR VPWR fd._1013_ sky130_fd_sc_hd__mux2_1
XFILLER_161_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._7635_ fd._2743_ fd._2924_ fd._2874_ VGND VGND VPWR VPWR fd._2926_ sky130_fd_sc_hd__mux2_1
XFILLER_12_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4847_ fd._3936_ fd._3940_ VGND VGND VPWR VPWR fd._3941_ sky130_fd_sc_hd__xnor2_1
XFILLER_115_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_150 VGND VGND VPWR VPWR user_project_wrapper_150/HI la_data_out[28]
+ sky130_fd_sc_hd__conb_1
XFILLER_177_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_project_wrapper_161 VGND VGND VPWR VPWR user_project_wrapper_161/HI la_data_out[39]
+ sky130_fd_sc_hd__conb_1
Xuser_project_wrapper_172 VGND VGND VPWR VPWR user_project_wrapper_172/HI la_data_out[50]
+ sky130_fd_sc_hd__conb_1
XFILLER_82_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._7566_ fd._2849_ VGND VGND VPWR VPWR fd._2850_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_115_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_183 VGND VGND VPWR VPWR user_project_wrapper_183/HI la_data_out[61]
+ sky130_fd_sc_hd__conb_1
Xfd._4778_ fd._3696_ fd._3871_ VGND VGND VPWR VPWR fd._3872_ sky130_fd_sc_hd__xnor2_1
XFILLER_173_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_194 VGND VGND VPWR VPWR user_project_wrapper_194/HI la_data_out[72]
+ sky130_fd_sc_hd__conb_1
XFILLER_86_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6517_ fd._1691_ fd._1695_ fd._1615_ VGND VGND VPWR VPWR fd._1696_ sky130_fd_sc_hd__mux2_1
XFILLER_141_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7497_ fd._2538_ fd._2561_ VGND VGND VPWR VPWR fd._2774_ sky130_fd_sc_hd__and2_1
XFILLER_87_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6448_ fd._1505_ fd._1619_ VGND VGND VPWR VPWR fd._1620_ sky130_fd_sc_hd__xnor2_1
XFILLER_25_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6379_ fd._1377_ fd._1404_ VGND VGND VPWR VPWR fd._1544_ sky130_fd_sc_hd__nand2_1
XFILLER_95_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8118_ fd.b\[24\] fd.a\[24\] VGND VGND VPWR VPWR fd._3433_ sky130_fd_sc_hd__and2b_1
XFILLER_186_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_270_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_266_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8049_ fd._1286_ fd._3380_ fd._3374_ fd._2427_ VGND VGND VPWR VPWR fd._3381_ sky130_fd_sc_hd__a22oi_1
XFILLER_270_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_260_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_9149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_1591 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_273_1556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_267_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput15 io_in[22] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_4
XFILLER_7_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput26 io_in[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_4
XFILLER_183_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5750_ fd._0771_ VGND VGND VPWR VPWR fd._0852_ sky130_fd_sc_hd__inv_2
XFILLER_7_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4701_ fd._3035_ fd._3794_ VGND VGND VPWR VPWR fd._3795_ sky130_fd_sc_hd__or2_1
Xfd._5681_ fd._0479_ fd._0774_ VGND VGND VPWR VPWR fd._0776_ sky130_fd_sc_hd__or2_1
XFILLER_100_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_8960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7420_ fd._1645_ fd._2608_ VGND VGND VPWR VPWR fd._2689_ sky130_fd_sc_hd__xnor2_1
XTAP_8971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4632_ fd._3557_ fd._3725_ VGND VGND VPWR VPWR fd._3726_ sky130_fd_sc_hd__xor2_1
XTAP_8982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._7351_ fd._2076_ fd._2612_ VGND VGND VPWR VPWR fd._2613_ sky130_fd_sc_hd__xnor2_1
XFILLER_123_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_257_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4563_ fd._3510_ fd._3656_ fd._3508_ VGND VGND VPWR VPWR fd._3657_ sky130_fd_sc_hd__o21ai_1
XFILLER_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6302_ fd._1456_ fd._1457_ fd._1458_ fd._1454_ VGND VGND VPWR VPWR fd._1459_ sky130_fd_sc_hd__a31o_1
XFILLER_250_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7282_ fd._2366_ fd._2536_ fd._2505_ VGND VGND VPWR VPWR fd._2537_ sky130_fd_sc_hd__mux2_1
Xfd._4494_ fd.b\[19\] fd._3587_ VGND VGND VPWR VPWR fd._3588_ sky130_fd_sc_hd__nand2_1
XFILLER_270_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6233_ fd._0450_ fd._1382_ VGND VGND VPWR VPWR fd._1383_ sky130_fd_sc_hd__or2_1
XFILLER_265_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_226_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6164_ fd._1304_ fd._1306_ VGND VGND VPWR VPWR fd._1307_ sky130_fd_sc_hd__nor2_1
XFILLER_77_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_281_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5115_ fd._3905_ fd._0152_ VGND VGND VPWR VPWR fd._0154_ sky130_fd_sc_hd__or2_1
XFILLER_111_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_279_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6095_ fd._1223_ VGND VGND VPWR VPWR fd._1232_ sky130_fd_sc_hd__buf_6
XFILLER_209_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5046_ fd._4035_ fd._0077_ VGND VGND VPWR VPWR fd._0078_ sky130_fd_sc_hd__xnor2_1
XFILLER_221_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6997_ fd._2093_ fd._2117_ VGND VGND VPWR VPWR fd._2224_ sky130_fd_sc_hd__nand2_1
XFILLER_146_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5948_ fd._2738_ fd._1051_ VGND VGND VPWR VPWR fd._1070_ sky130_fd_sc_hd__or2_1
XFILLER_228_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5879_ fd._0991_ fd._0993_ VGND VGND VPWR VPWR fd._0994_ sky130_fd_sc_hd__xor2_1
XFILLER_161_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_255_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1690 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._7618_ fd._2326_ fd._2905_ VGND VGND VPWR VPWR fd._2907_ sky130_fd_sc_hd__and2_1
XFILLER_192_1554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7549_ fd._2640_ VGND VGND VPWR VPWR fd._2831_ sky130_fd_sc_hd__clkinv_2
XFILLER_276_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_284_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_243_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_249_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_1410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_273_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_8278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_279_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_281_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_263_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_267_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_1444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6920_ fd._2136_ fd._2138_ fd._2116_ VGND VGND VPWR VPWR fd._2139_ sky130_fd_sc_hd__mux2_1
XFILLER_124_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6851_ fd._2054_ fd._2062_ VGND VGND VPWR VPWR fd._2063_ sky130_fd_sc_hd__nor2_1
XFILLER_129_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5802_ fd._0662_ fd._0908_ VGND VGND VPWR VPWR fd._0909_ sky130_fd_sc_hd__nor2_1
XFILLER_184_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_229_ fd.c\[21\] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_1
XFILLER_129_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6782_ fd._1750_ fd._1776_ fd._1746_ VGND VGND VPWR VPWR fd._1987_ sky130_fd_sc_hd__o21a_1
XFILLER_176_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5733_ fd._0638_ fd._0830_ fd._0832_ VGND VGND VPWR VPWR fd._0833_ sky130_fd_sc_hd__o21bai_1
XFILLER_195_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5664_ fd._0592_ fd._0599_ VGND VGND VPWR VPWR fd._0757_ sky130_fd_sc_hd__xnor2_1
XFILLER_170_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_256_1584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._4615_ fd._3708_ fd._3704_ VGND VGND VPWR VPWR fd._3709_ sky130_fd_sc_hd__and2_1
XFILLER_252_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7403_ fd._2629_ fd._2659_ fd._2669_ VGND VGND VPWR VPWR fd._2670_ sky130_fd_sc_hd__a21o_2
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5595_ fd._1341_ fd._0680_ VGND VGND VPWR VPWR fd._0682_ sky130_fd_sc_hd__xnor2_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7334_ fd._2593_ VGND VGND VPWR VPWR fd._2594_ sky130_fd_sc_hd__inv_2
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4546_ fd._3638_ fd._3639_ fd._3422_ VGND VGND VPWR VPWR fd._3640_ sky130_fd_sc_hd__a21boi_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_273_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7265_ fd._2388_ fd._2355_ VGND VGND VPWR VPWR fd._2519_ sky130_fd_sc_hd__and2b_1
XFILLER_22_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4477_ fd._2617_ fd._3570_ fd._3211_ VGND VGND VPWR VPWR fd._3571_ sky130_fd_sc_hd__mux2_1
XFILLER_214_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6216_ fd._0807_ fd._1188_ VGND VGND VPWR VPWR fd._1365_ sky130_fd_sc_hd__or2_1
XFILLER_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7196_ fd._2266_ fd._2442_ fd._2323_ VGND VGND VPWR VPWR fd._2443_ sky130_fd_sc_hd__mux2_1
XFILLER_25_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_285_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6147_ fd._1319_ fd._1288_ VGND VGND VPWR VPWR fd._1289_ sky130_fd_sc_hd__or2_1
XFILLER_80_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_253_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6078_ fd._0821_ fd._1210_ fd._1204_ fd._0318_ fd._1212_ VGND VGND VPWR VPWR fd._1213_
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5029_ fd._0058_ VGND VGND VPWR VPWR fd._0059_ sky130_fd_sc_hd__buf_6
XFILLER_221_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_257_1359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_270_1515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_276_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_268_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_271_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_260_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_1639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4400_ fd._3491_ fd._3493_ VGND VGND VPWR VPWR fd._3494_ sky130_fd_sc_hd__xnor2_1
XFILLER_239_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5380_ fd._4011_ fd._0444_ fd._0442_ fd._0125_ VGND VGND VPWR VPWR fd._0445_ sky130_fd_sc_hd__o22ai_1
XTAP_6673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4331_ fd._1363_ fd._0978_ VGND VGND VPWR VPWR fd._2826_ sky130_fd_sc_hd__nor2_1
XFILLER_255_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7050_ fd._2279_ fd._2281_ VGND VGND VPWR VPWR fd._2282_ sky130_fd_sc_hd__xnor2_1
Xfd._4262_ fd.b\[6\] fd._1693_ VGND VGND VPWR VPWR fd._2067_ sky130_fd_sc_hd__nor2_1
XFILLER_212_1498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6001_ fd._4055_ fd._0957_ VGND VGND VPWR VPWR fd._1128_ sky130_fd_sc_hd__xnor2_1
XFILLER_223_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4193_ fd._1297_ VGND VGND VPWR VPWR fd._1308_ sky130_fd_sc_hd__buf_6
XFILLER_21_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_250_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7952_ fd._2377_ fd._3170_ VGND VGND VPWR VPWR fd._3274_ sky130_fd_sc_hd__or2_1
XFILLER_31_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6903_ fd._2005_ fd._2118_ VGND VGND VPWR VPWR fd._2120_ sky130_fd_sc_hd__or2_1
XFILLER_15_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7883_ fd._1661_ fd._3115_ VGND VGND VPWR VPWR fd._3198_ sky130_fd_sc_hd__nor2_1
XFILLER_129_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6834_ fd._2037_ fd._2042_ fd._2043_ VGND VGND VPWR VPWR fd._2044_ sky130_fd_sc_hd__a21o_1
XFILLER_239_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6765_ fd._1967_ VGND VGND VPWR VPWR fd._1969_ sky130_fd_sc_hd__buf_6
XFILLER_128_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5716_ fd._0811_ fd._0814_ VGND VGND VPWR VPWR fd._0815_ sky130_fd_sc_hd__xor2_1
XFILLER_239_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6696_ fd._1668_ fd._1673_ VGND VGND VPWR VPWR fd._1893_ sky130_fd_sc_hd__xnor2_1
XFILLER_131_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_258_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5647_ fd._0731_ fd._0737_ fd._0738_ VGND VGND VPWR VPWR fd._0739_ sky130_fd_sc_hd__a21o_1
XFILLER_131_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5578_ fd._0533_ fd._0531_ VGND VGND VPWR VPWR fd._0663_ sky130_fd_sc_hd__nand2_1
XFILLER_135_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4529_ fd._3604_ fd._3618_ fd._3619_ fd._3622_ VGND VGND VPWR VPWR fd._3623_ sky130_fd_sc_hd__a31o_1
Xfd._7317_ fd._2517_ fd._2523_ fd._2565_ fd._2574_ fd._2575_ VGND VGND VPWR VPWR fd._2576_
+ sky130_fd_sc_hd__a41o_1
XFILLER_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_285_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7248_ fd._2494_ fd._2487_ fd._2499_ VGND VGND VPWR VPWR fd._2500_ sky130_fd_sc_hd__o21ai_1
XFILLER_2_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_253_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7179_ fd._2255_ fd._2422_ fd._2423_ VGND VGND VPWR VPWR fd._2424_ sky130_fd_sc_hd__mux2_1
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_257_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_268_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_277_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4880_ fd._3897_ fd._3973_ VGND VGND VPWR VPWR fd._3974_ sky130_fd_sc_hd__xnor2_1
XFILLER_201_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_279_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6550_ fd._1731_ VGND VGND VPWR VPWR fd._1732_ sky130_fd_sc_hd__inv_2
XFILLER_99_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5501_ fd._1308_ fd._0576_ VGND VGND VPWR VPWR fd._0578_ sky130_fd_sc_hd__and2_1
XFILLER_253_1543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6481_ fd._0846_ VGND VGND VPWR VPWR fd._1656_ sky130_fd_sc_hd__buf_6
XFILLER_113_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8220_ net73 net4 VGND VGND VPWR VPWR fd.a\[12\] sky130_fd_sc_hd__dfxtp_1
Xfd._5432_ fd._0089_ fd._0495_ VGND VGND VPWR VPWR fd._0502_ sky130_fd_sc_hd__and2_1
XTAP_7193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8151_ fd._3456_ fd._3465_ VGND VGND VPWR VPWR fd._3466_ sky130_fd_sc_hd__nand2_1
XTAP_6492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5363_ fd._0251_ fd._0266_ fd._0425_ VGND VGND VPWR VPWR fd._0426_ sky130_fd_sc_hd__mux2_1
XFILLER_209_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7102_ fd._1600_ fd._2338_ VGND VGND VPWR VPWR fd._2339_ sky130_fd_sc_hd__or2_1
XFILLER_282_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4314_ fd._2584_ fd._2628_ VGND VGND VPWR VPWR fd._2639_ sky130_fd_sc_hd__or2_1
XFILLER_255_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8082_ fd._1813_ fd._2020_ fd._3398_ VGND VGND VPWR VPWR fd._3408_ sky130_fd_sc_hd__mux2_1
XFILLER_76_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5294_ fd._0303_ fd._0342_ fd._0348_ fd._0349_ VGND VGND VPWR VPWR fd._0350_ sky130_fd_sc_hd__a31o_1
XFILLER_3_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._7033_ fd._2262_ fd._2088_ VGND VGND VPWR VPWR fd._2263_ sky130_fd_sc_hd__nor2_1
Xfd._4245_ fd._1858_ fd._1869_ fd._1209_ VGND VGND VPWR VPWR fd._1880_ sky130_fd_sc_hd__mux2_1
XFILLER_235_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_251_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4176_ fd._1110_ VGND VGND VPWR VPWR fd._1121_ sky130_fd_sc_hd__clkinv_4
XFILLER_264_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_251_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_1656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7935_ fd._3249_ fd._3253_ fd._3254_ VGND VGND VPWR VPWR fd._3256_ sky130_fd_sc_hd__and3_1
XFILLER_143_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7866_ fd._3149_ fd._3152_ fd._3177_ fd._3179_ fd._3147_ VGND VGND VPWR VPWR fd._3180_
+ sky130_fd_sc_hd__o311a_1
XFILLER_258_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1700 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6817_ fd._1816_ fd._2025_ VGND VGND VPWR VPWR fd._2026_ sky130_fd_sc_hd__nor2_1
XFILLER_145_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7797_ fd._1330_ fd._3098_ VGND VGND VPWR VPWR fd._3104_ sky130_fd_sc_hd__and2_1
XFILLER_236_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._6748_ fd._1761_ VGND VGND VPWR VPWR fd._1950_ sky130_fd_sc_hd__clkinv_2
XFILLER_160_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6679_ fd._1650_ fd._1873_ VGND VGND VPWR VPWR fd._1874_ sky130_fd_sc_hd__nand2_1
XFILLER_132_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_274_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_219_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_276_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_272_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_264_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5981_ fd._0941_ fd._0939_ VGND VGND VPWR VPWR fd._1106_ sky130_fd_sc_hd__nor2_1
XFILLER_119_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7720_ fd._2887_ fd._2893_ fd._3018_ fd._2885_ VGND VGND VPWR VPWR fd._3019_ sky130_fd_sc_hd__o31ai_1
Xfd._4932_ fd._3708_ fd._4023_ VGND VGND VPWR VPWR fd._4026_ sky130_fd_sc_hd__and2_1
XFILLER_145_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4863_ fd._3956_ fd._3955_ fd._3763_ VGND VGND VPWR VPWR fd._3957_ sky130_fd_sc_hd__mux2_1
XFILLER_145_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7651_ fd._1751_ fd._2941_ VGND VGND VPWR VPWR fd._2943_ sky130_fd_sc_hd__nand2_1
XFILLER_127_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6602_ fd._1602_ VGND VGND VPWR VPWR fd._1789_ sky130_fd_sc_hd__clkinv_2
XFILLER_142_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4794_ fd._3858_ fd._3862_ fd._3885_ fd._3887_ VGND VGND VPWR VPWR fd._3888_ sky130_fd_sc_hd__a31o_1
Xfd._7582_ fd._2845_ fd._2836_ fd._2844_ VGND VGND VPWR VPWR fd._2867_ sky130_fd_sc_hd__a21oi_1
XFILLER_114_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6533_ fd._1642_ VGND VGND VPWR VPWR fd._1713_ sky130_fd_sc_hd__inv_2
XFILLER_114_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6464_ fd._1632_ fd._1636_ VGND VGND VPWR VPWR fd._1637_ sky130_fd_sc_hd__nand2_1
XFILLER_151_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5415_ fd._0295_ VGND VGND VPWR VPWR fd._0484_ sky130_fd_sc_hd__clkinv_2
XFILLER_214_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._8203_ net68 fd.ec\[4\] VGND VGND VPWR VPWR fd.c\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6395_ fd._1402_ fd._1383_ VGND VGND VPWR VPWR fd._1562_ sky130_fd_sc_hd__or2b_1
XFILLER_95_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8134_ fd._3447_ fd._3448_ VGND VGND VPWR VPWR fd.ec\[2\] sky130_fd_sc_hd__nand2_1
Xfd._5346_ fd._0069_ fd._0407_ fd._0270_ VGND VGND VPWR VPWR fd._0408_ sky130_fd_sc_hd__mux2_1
XFILLER_55_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8065_ fd._3189_ VGND VGND VPWR VPWR fd._3398_ sky130_fd_sc_hd__buf_6
XFILLER_236_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5277_ fd._0100_ fd._0331_ VGND VGND VPWR VPWR fd._0332_ sky130_fd_sc_hd__nand2_1
XFILLER_222_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_282_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4228_ fd._1638_ fd._1682_ fd._1209_ VGND VGND VPWR VPWR fd._1693_ sky130_fd_sc_hd__mux2_1
XFILLER_212_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7016_ fd._1816_ fd._2244_ VGND VGND VPWR VPWR fd._2245_ sky130_fd_sc_hd__nor2_1
XFILLER_149_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4159_ fd._0725_ fd._0769_ fd._0923_ VGND VGND VPWR VPWR fd._0934_ sky130_fd_sc_hd__or3_1
XFILLER_260_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7918_ fd._3236_ fd._3232_ fd._3077_ fd._3036_ VGND VGND VPWR VPWR fd._3237_ sky130_fd_sc_hd__o211a_1
XFILLER_17_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7849_ fd._2959_ fd._3160_ VGND VGND VPWR VPWR fd._3161_ sky130_fd_sc_hd__xnor2_1
XTAP_8619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_1530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_273_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_258_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_1560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_261_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_261_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_243_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_272_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5200_ fd._0246_ VGND VGND VPWR VPWR fd._0247_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_92_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6180_ fd._1162_ fd._1324_ fd._1232_ VGND VGND VPWR VPWR fd._1325_ sky130_fd_sc_hd__nand3_1
XTAP_4150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5131_ fd._0169_ fd._0170_ fd._0060_ VGND VGND VPWR VPWR fd._0171_ sky130_fd_sc_hd__a21o_1
XFILLER_168_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_264_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5062_ fd._0093_ fd._0094_ VGND VGND VPWR VPWR fd._0095_ sky130_fd_sc_hd__xnor2_1
XFILLER_61_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_1607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_261_1620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5964_ fd._0662_ fd._1086_ VGND VGND VPWR VPWR fd._1087_ sky130_fd_sc_hd__nor2_1
XFILLER_146_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7703_ fd._1645_ fd._2697_ VGND VGND VPWR VPWR fd._3000_ sky130_fd_sc_hd__and2_1
Xfd._4915_ fd._3954_ fd._3958_ fd._4007_ fd._4008_ VGND VGND VPWR VPWR fd._4009_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_174_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5895_ fd._1008_ fd._1010_ VGND VGND VPWR VPWR fd._1012_ sky130_fd_sc_hd__xor2_1
XFILLER_179_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7634_ fd._2921_ fd._2923_ VGND VGND VPWR VPWR fd._2924_ sky130_fd_sc_hd__xnor2_1
XFILLER_127_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._4846_ fd._3938_ fd._3939_ VGND VGND VPWR VPWR fd._3940_ sky130_fd_sc_hd__nor2_1
XFILLER_115_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_project_wrapper_140 VGND VGND VPWR VPWR user_project_wrapper_140/HI la_data_out[18]
+ sky130_fd_sc_hd__conb_1
XFILLER_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_255_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xuser_project_wrapper_151 VGND VGND VPWR VPWR user_project_wrapper_151/HI la_data_out[29]
+ sky130_fd_sc_hd__conb_1
XFILLER_217_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_162 VGND VGND VPWR VPWR user_project_wrapper_162/HI la_data_out[40]
+ sky130_fd_sc_hd__conb_1
XFILLER_255_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_project_wrapper_173 VGND VGND VPWR VPWR user_project_wrapper_173/HI la_data_out[51]
+ sky130_fd_sc_hd__conb_1
XFILLER_255_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7565_ fd._2465_ fd._2828_ VGND VGND VPWR VPWR fd._2849_ sky130_fd_sc_hd__and2_1
Xfd._4777_ fd._3870_ fd._3694_ VGND VGND VPWR VPWR fd._3871_ sky130_fd_sc_hd__nand2_1
XFILLER_115_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_184 VGND VGND VPWR VPWR user_project_wrapper_184/HI la_data_out[62]
+ sky130_fd_sc_hd__conb_1
XFILLER_82_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_project_wrapper_195 VGND VGND VPWR VPWR user_project_wrapper_195/HI la_data_out[73]
+ sky130_fd_sc_hd__conb_1
XFILLER_173_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6516_ fd._1493_ fd._1694_ VGND VGND VPWR VPWR fd._1695_ sky130_fd_sc_hd__nand2_1
XFILLER_130_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7496_ fd._2737_ fd._2742_ fd._2770_ fd._2772_ VGND VGND VPWR VPWR fd._2773_ sky130_fd_sc_hd__a31o_1
XFILLER_25_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6447_ fd._1512_ fd._1511_ VGND VGND VPWR VPWR fd._1619_ sky130_fd_sc_hd__and2b_1
XFILLER_151_1444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6378_ fd._1541_ fd._1542_ VGND VGND VPWR VPWR fd._1543_ sky130_fd_sc_hd__and2_1
XFILLER_55_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8117_ fd.a\[24\] fd.b\[24\] VGND VGND VPWR VPWR fd._3432_ sky130_fd_sc_hd__and2b_1
XFILLER_244_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5329_ fd._1264_ fd._0073_ VGND VGND VPWR VPWR fd._0389_ sky130_fd_sc_hd__nand2_1
XFILLER_110_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8048_ fd._3207_ fd._3241_ fd._3377_ fd._3379_ VGND VGND VPWR VPWR fd._3380_ sky130_fd_sc_hd__a31oi_1
XFILLER_110_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_270_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_266_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_252_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_260_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_273_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_262_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput16 io_in[23] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_1
XFILLER_128_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput27 io_in[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_4
XFILLER_11_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4700_ fd._3793_ fd._3627_ fd._3788_ VGND VGND VPWR VPWR fd._3794_ sky130_fd_sc_hd__mux2_1
XFILLER_202_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5680_ fd._0479_ fd._0774_ VGND VGND VPWR VPWR fd._0775_ sky130_fd_sc_hd__nand2_1
XFILLER_183_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4631_ fd._3555_ fd._3724_ fd._3625_ VGND VGND VPWR VPWR fd._3725_ sky130_fd_sc_hd__nand3_1
XFILLER_269_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_8994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4562_ fd._3514_ fd._3543_ VGND VGND VPWR VPWR fd._3656_ sky130_fd_sc_hd__or2_1
Xfd._7350_ fd._2610_ fd._2577_ fd._2611_ VGND VGND VPWR VPWR fd._2612_ sky130_fd_sc_hd__o21a_1
XFILLER_112_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6301_ fd._1405_ fd._1411_ fd._1417_ fd._1412_ fd._1361_ VGND VGND VPWR VPWR fd._1458_
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_61_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7281_ fd._2534_ fd._2535_ VGND VGND VPWR VPWR fd._2536_ sky130_fd_sc_hd__xnor2_1
Xfd._4493_ fd._2936_ fd._3586_ fd._3222_ VGND VGND VPWR VPWR fd._3587_ sky130_fd_sc_hd__mux2_1
XFILLER_84_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6232_ fd._1204_ fd._1381_ fd._1349_ VGND VGND VPWR VPWR fd._1382_ sky130_fd_sc_hd__mux2_1
XFILLER_38_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6163_ fd._1159_ fd._1305_ fd._1232_ VGND VGND VPWR VPWR fd._1306_ sky130_fd_sc_hd__mux2_1
XFILLER_19_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5114_ fd._0151_ fd._3975_ fd._0060_ VGND VGND VPWR VPWR fd._0152_ sky130_fd_sc_hd__mux2_1
XFILLER_168_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6094_ fd._1140_ fd._1147_ VGND VGND VPWR VPWR fd._1230_ sky130_fd_sc_hd__xor2_1
XTAP_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5045_ fd._4041_ fd._4039_ VGND VGND VPWR VPWR fd._0077_ sky130_fd_sc_hd__and2b_1
XFILLER_209_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6996_ fd._2093_ fd._2117_ VGND VGND VPWR VPWR fd._2223_ sky130_fd_sc_hd__or2_1
XFILLER_179_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5947_ fd._1088_ fd._1068_ VGND VGND VPWR VPWR fd._1069_ sky130_fd_sc_hd__and2_1
XFILLER_105_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5878_ fd._0810_ fd._0992_ VGND VGND VPWR VPWR fd._0993_ sky130_fd_sc_hd__nand2_1
XFILLER_259_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7617_ fd._2326_ fd._2905_ VGND VGND VPWR VPWR fd._2906_ sky130_fd_sc_hd__nor2_1
XFILLER_115_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4829_ fd._3823_ fd._3828_ fd._3922_ VGND VGND VPWR VPWR fd._3923_ sky130_fd_sc_hd__or3_1
XFILLER_216_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7548_ fd._2829_ VGND VGND VPWR VPWR fd._2830_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_244_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_276_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_275_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7479_ fd._0821_ fd._2556_ VGND VGND VPWR VPWR fd._2754_ sky130_fd_sc_hd__xnor2_1
XTAP_4919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_262_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_285_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_256_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_1439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_273_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_267_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_249_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._6850_ fd._1304_ fd._2052_ fd._2061_ fd._1431_ VGND VGND VPWR VPWR fd._2062_ sky130_fd_sc_hd__o22a_1
XFILLER_50_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_228_ fd.c\[20\] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_1
Xfd._5801_ fd._0675_ fd._0907_ fd._0801_ VGND VGND VPWR VPWR fd._0908_ sky130_fd_sc_hd__mux2_1
XFILLER_200_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6781_ fd._1943_ fd._1949_ fd._1985_ fd._1941_ VGND VGND VPWR VPWR fd._1986_ sky130_fd_sc_hd__o31a_1
XFILLER_129_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5732_ fd._3537_ fd._0829_ VGND VGND VPWR VPWR fd._0832_ sky130_fd_sc_hd__and2_1
XFILLER_7_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_256_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5663_ fd._0653_ fd._0749_ fd._0753_ fd._0594_ VGND VGND VPWR VPWR fd._0756_ sky130_fd_sc_hd__a31o_1
XFILLER_139_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7402_ fd._2665_ fd._2668_ VGND VGND VPWR VPWR fd._2669_ sky130_fd_sc_hd__or2b_1
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4614_ fd._0428_ VGND VGND VPWR VPWR fd._3708_ sky130_fd_sc_hd__buf_6
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5594_ fd._0519_ fd._0679_ fd._0614_ VGND VGND VPWR VPWR fd._0680_ sky130_fd_sc_hd__mux2_1
XFILLER_174_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7333_ fd._2591_ fd._2592_ VGND VGND VPWR VPWR fd._2593_ sky130_fd_sc_hd__and2_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4545_ fd._3560_ VGND VGND VPWR VPWR fd._3639_ sky130_fd_sc_hd__inv_2
XFILLER_257_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4476_ fd._2573_ fd._2661_ VGND VGND VPWR VPWR fd._3570_ sky130_fd_sc_hd__xnor2_1
Xfd._7264_ fd._2515_ fd._2516_ VGND VGND VPWR VPWR fd._2517_ sky130_fd_sc_hd__nor2_1
XFILLER_226_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6215_ fd._1196_ fd._1205_ fd._1213_ fd._1214_ VGND VGND VPWR VPWR fd._1364_ sky130_fd_sc_hd__a31o_1
XFILLER_281_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7195_ fd._2440_ fd._2269_ VGND VGND VPWR VPWR fd._2442_ sky130_fd_sc_hd__xnor2_1
XFILLER_93_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_285_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_281_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6146_ fd._1284_ fd._1223_ fd._1287_ VGND VGND VPWR VPWR fd._1288_ sky130_fd_sc_hd__a21oi_1
XFILLER_267_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6077_ fd._0821_ fd._1208_ fd._1206_ fd._1211_ VGND VGND VPWR VPWR fd._1212_ sky130_fd_sc_hd__o211a_1
XFILLER_263_1556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5028_ fd._0050_ fd._0052_ fd._0057_ VGND VGND VPWR VPWR fd._0058_ sky130_fd_sc_hd__and3_1
XFILLER_228_1698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_279_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6979_ fd._2203_ VGND VGND VPWR VPWR fd._2204_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_146_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_276_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_271_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_268_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_260_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_271_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_281_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_279_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4330_ fd.a\[19\] VGND VGND VPWR VPWR fd._2815_ sky130_fd_sc_hd__clkinv_2
XTAP_6696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_251_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4261_ fd._1847_ fd._2023_ fd._2034_ fd._2045_ VGND VGND VPWR VPWR fd._2056_ sky130_fd_sc_hd__a211o_1
XFILLER_247_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_282_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6000_ fd._1117_ fd._1125_ fd._1126_ VGND VGND VPWR VPWR fd._1127_ sky130_fd_sc_hd__o21ba_1
XFILLER_262_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_263_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4192_ fd.b\[15\] VGND VGND VPWR VPWR fd._1297_ sky130_fd_sc_hd__buf_6
XFILLER_207_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7951_ fd._3171_ fd._3272_ VGND VGND VPWR VPWR fd._3273_ sky130_fd_sc_hd__xnor2_1
XFILLER_128_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6902_ fd._2005_ fd._2118_ VGND VGND VPWR VPWR fd._2119_ sky130_fd_sc_hd__nand2_1
XFILLER_30_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7882_ fd._1797_ fd._3128_ fd._3190_ fd._3195_ fd._3196_ VGND VGND VPWR VPWR fd._3197_
+ sky130_fd_sc_hd__a221o_1
XFILLER_276_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6833_ fd._1242_ fd._2036_ VGND VGND VPWR VPWR fd._2043_ sky130_fd_sc_hd__nor2_1
XFILLER_129_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_278_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6764_ fd._1821_ fd._1835_ fd._1915_ VGND VGND VPWR VPWR fd._1967_ sky130_fd_sc_hd__and3_1
XFILLER_143_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5715_ fd._0630_ fd._0812_ VGND VGND VPWR VPWR fd._0814_ sky130_fd_sc_hd__nand2_1
Xfd._6695_ fd._1871_ fd._1886_ fd._1890_ VGND VGND VPWR VPWR fd._1892_ sky130_fd_sc_hd__a21oi_1
XFILLER_131_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5646_ fd._1308_ fd._0735_ VGND VGND VPWR VPWR fd._0738_ sky130_fd_sc_hd__and2_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5577_ fd._3980_ VGND VGND VPWR VPWR fd._0662_ sky130_fd_sc_hd__buf_6
XFILLER_154_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7316_ fd._2572_ fd._2515_ fd._2571_ VGND VGND VPWR VPWR fd._2575_ sky130_fd_sc_hd__o21ba_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4528_ fd._3611_ fd._3617_ fd._3620_ fd._3621_ VGND VGND VPWR VPWR fd._3622_ sky130_fd_sc_hd__o22ai_1
XFILLER_22_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7247_ fd._1242_ fd._2491_ VGND VGND VPWR VPWR fd._2499_ sky130_fd_sc_hd__or2_1
Xfd._4459_ fd._3498_ fd._3549_ fd._3552_ VGND VGND VPWR VPWR fd._3553_ sky130_fd_sc_hd__a21o_1
XFILLER_54_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_265_1607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7178_ fd._2323_ VGND VGND VPWR VPWR fd._2423_ sky130_fd_sc_hd__buf_6
XFILLER_0_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6129_ fd._1102_ fd._1100_ VGND VGND VPWR VPWR fd._1269_ sky130_fd_sc_hd__and2_1
XFILLER_55_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_263_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_257_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_270_1379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_268_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_260_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_1573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5500_ fd._1308_ fd._0576_ VGND VGND VPWR VPWR fd._0577_ sky130_fd_sc_hd__or2_1
XFILLER_153_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._6480_ fd._0846_ fd._1654_ VGND VGND VPWR VPWR fd._1655_ sky130_fd_sc_hd__nand2_1
XTAP_7161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._5431_ fd._3980_ fd._0500_ VGND VGND VPWR VPWR fd._0501_ sky130_fd_sc_hd__or2_1
XTAP_7183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8150_ fd._3463_ fd._3464_ VGND VGND VPWR VPWR fd._3465_ sky130_fd_sc_hd__or2_1
XTAP_6482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5362_ fd._0280_ fd._0413_ fd._0419_ fd._0424_ VGND VGND VPWR VPWR fd._0425_ sky130_fd_sc_hd__a31o_4
XTAP_6493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7101_ fd._2130_ fd._2337_ fd._2322_ VGND VGND VPWR VPWR fd._2338_ sky130_fd_sc_hd__mux2_1
XFILLER_3_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4313_ fd._2595_ fd._2617_ fd._1231_ VGND VGND VPWR VPWR fd._2628_ sky130_fd_sc_hd__mux2_1
XFILLER_208_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5293_ fd._0868_ fd._0347_ VGND VGND VPWR VPWR fd._0349_ sky130_fd_sc_hd__nor2_1
Xfd._8081_ fd._3407_ VGND VGND VPWR VPWR fd.mc\[8\] sky130_fd_sc_hd__clkbuf_1
XFILLER_23_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7032_ fd._2093_ fd._2087_ VGND VGND VPWR VPWR fd._2262_ sky130_fd_sc_hd__and2_1
Xfd._4244_ fd._0351_ fd._0395_ VGND VGND VPWR VPWR fd._1869_ sky130_fd_sc_hd__xnor2_1
XFILLER_224_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_250_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4175_ fd._0010_ fd._1099_ VGND VGND VPWR VPWR fd._1110_ sky130_fd_sc_hd__nor2_1
XFILLER_211_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_251_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_250_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_264_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7934_ fd._2863_ fd._3252_ VGND VGND VPWR VPWR fd._3254_ sky130_fd_sc_hd__nand2_1
XFILLER_52_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_223_1370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7865_ fd._2135_ fd._3139_ VGND VGND VPWR VPWR fd._3179_ sky130_fd_sc_hd__nand2_1
XFILLER_176_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6816_ fd._2022_ fd._2024_ fd._2020_ VGND VGND VPWR VPWR fd._2025_ sky130_fd_sc_hd__mux2_1
XFILLER_191_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7796_ fd._2076_ fd._3102_ VGND VGND VPWR VPWR fd._3103_ sky130_fd_sc_hd__or2_1
XFILLER_145_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6747_ fd._0312_ fd._1948_ VGND VGND VPWR VPWR fd._1949_ sky130_fd_sc_hd__nor2_1
XFILLER_219_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_271_1600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6678_ fd._1657_ fd._1655_ VGND VGND VPWR VPWR fd._1873_ sky130_fd_sc_hd__and2b_1
XFILLER_259_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5629_ fd._0718_ VGND VGND VPWR VPWR fd._0719_ sky130_fd_sc_hd__clkinv_4
XFILLER_131_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_1584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_227_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_1590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5980_ fd._0918_ fd._0935_ VGND VGND VPWR VPWR fd._1105_ sky130_fd_sc_hd__nand2_1
XFILLER_144_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_1519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._4931_ fd._3469_ fd._3975_ VGND VGND VPWR VPWR fd._4025_ sky130_fd_sc_hd__xnor2_1
XFILLER_201_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7650_ fd._1751_ fd._2941_ VGND VGND VPWR VPWR fd._2942_ sky130_fd_sc_hd__or2_1
Xfd._4862_ fd._3955_ fd._3800_ VGND VGND VPWR VPWR fd._3956_ sky130_fd_sc_hd__nand2_1
XFILLER_173_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6601_ fd._1732_ fd._1736_ fd._1778_ fd._1786_ fd._1787_ VGND VGND VPWR VPWR fd._1788_
+ sky130_fd_sc_hd__o41a_1
XFILLER_177_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7581_ fd._2856_ fd._2865_ VGND VGND VPWR VPWR fd._2866_ sky130_fd_sc_hd__and2_1
XFILLER_275_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4793_ fd._3886_ VGND VGND VPWR VPWR fd._3887_ sky130_fd_sc_hd__inv_2
XFILLER_153_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6532_ fd._1637_ fd._1710_ fd._1711_ VGND VGND VPWR VPWR fd._1712_ sky130_fd_sc_hd__and3_1
XFILLER_99_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._6463_ fd._1428_ fd._1617_ fd._1635_ VGND VGND VPWR VPWR fd._1636_ sky130_fd_sc_hd__o21a_1
XFILLER_113_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8202_ net66 fd.ec\[3\] VGND VGND VPWR VPWR fd.c\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_171_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5414_ fd._1352_ VGND VGND VPWR VPWR fd._0482_ sky130_fd_sc_hd__buf_6
XFILLER_151_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._6394_ fd._1382_ VGND VGND VPWR VPWR fd._1560_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_7_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_282_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8133_ fd._3436_ fd._3446_ VGND VGND VPWR VPWR fd._3448_ sky130_fd_sc_hd__or2_1
XFILLER_231_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._5345_ fd._0403_ fd._0405_ VGND VGND VPWR VPWR fd._0407_ sky130_fd_sc_hd__xnor2_1
XFILLER_209_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8064_ fd._3396_ VGND VGND VPWR VPWR fd.mc\[0\] sky130_fd_sc_hd__buf_4
Xfd._5276_ fd._0105_ fd._0135_ VGND VGND VPWR VPWR fd._0331_ sky130_fd_sc_hd__and2_1
XFILLER_184_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7015_ fd._2238_ fd._2240_ fd._2241_ fd._2242_ VGND VGND VPWR VPWR fd._2244_ sky130_fd_sc_hd__a31o_1
Xfd._4227_ fd._0274_ fd._1671_ VGND VGND VPWR VPWR fd._1682_ sky130_fd_sc_hd__xnor2_1
XFILLER_251_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1590 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4158_ fd._0747_ fd._0791_ VGND VGND VPWR VPWR fd._0923_ sky130_fd_sc_hd__nor2_1
XFILLER_71_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4089_ fd._0131_ fd.a\[19\] VGND VGND VPWR VPWR fd._0164_ sky130_fd_sc_hd__nor2_1
XFILLER_71_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7917_ fd._3034_ VGND VGND VPWR VPWR fd._3236_ sky130_fd_sc_hd__inv_2
XFILLER_192_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7848_ fd._3159_ fd._2957_ VGND VGND VPWR VPWR fd._3160_ sky130_fd_sc_hd__nor2_1
XTAP_8609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_254_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7779_ fd._3082_ fd._3083_ VGND VGND VPWR VPWR fd._3084_ sky130_fd_sc_hd__xnor2_1
XFILLER_69_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_258_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_259_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_273_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_261_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_265_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_243_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_276_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_269_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_285_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_264_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_280_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5130_ fd._4042_ fd._4046_ VGND VGND VPWR VPWR fd._0170_ sky130_fd_sc_hd__or2_1
XTAP_4173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5061_ fd._3993_ fd._4016_ VGND VGND VPWR VPWR fd._0094_ sky130_fd_sc_hd__and2b_1
XFILLER_233_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_261_1643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5963_ fd._0924_ fd._1085_ fd._0998_ VGND VGND VPWR VPWR fd._1086_ sky130_fd_sc_hd__mux2_1
XFILLER_179_1504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7702_ fd._2703_ fd._2801_ VGND VGND VPWR VPWR fd._2999_ sky130_fd_sc_hd__nand2_1
Xfd._4914_ fd._4001_ VGND VGND VPWR VPWR fd._4008_ sky130_fd_sc_hd__clkinv_2
XFILLER_179_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5894_ fd._1009_ fd._0834_ VGND VGND VPWR VPWR fd._1010_ sky130_fd_sc_hd__nor2_1
XFILLER_63_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7633_ fd._2742_ fd._2922_ VGND VGND VPWR VPWR fd._2923_ sky130_fd_sc_hd__nand2_1
Xfd._4845_ fd._3773_ fd._3789_ VGND VGND VPWR VPWR fd._3939_ sky130_fd_sc_hd__and2_1
XFILLER_161_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_130 VGND VGND VPWR VPWR user_project_wrapper_130/HI la_data_out[8]
+ sky130_fd_sc_hd__conb_1
XFILLER_154_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_project_wrapper_141 VGND VGND VPWR VPWR user_project_wrapper_141/HI la_data_out[19]
+ sky130_fd_sc_hd__conb_1
Xuser_project_wrapper_152 VGND VGND VPWR VPWR user_project_wrapper_152/HI la_data_out[30]
+ sky130_fd_sc_hd__conb_1
Xfd._7564_ fd._2839_ fd._2846_ VGND VGND VPWR VPWR fd._2847_ sky130_fd_sc_hd__and2_1
Xuser_project_wrapper_163 VGND VGND VPWR VPWR user_project_wrapper_163/HI la_data_out[41]
+ sky130_fd_sc_hd__conb_1
Xfd._4776_ fd._3688_ fd._3693_ VGND VGND VPWR VPWR fd._3870_ sky130_fd_sc_hd__or2_1
XFILLER_114_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_174 VGND VGND VPWR VPWR user_project_wrapper_174/HI la_data_out[52]
+ sky130_fd_sc_hd__conb_1
XFILLER_130_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_185 VGND VGND VPWR VPWR user_project_wrapper_185/HI la_data_out[63]
+ sky130_fd_sc_hd__conb_1
XFILLER_233_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_project_wrapper_196 VGND VGND VPWR VPWR user_project_wrapper_196/HI la_data_out[74]
+ sky130_fd_sc_hd__conb_1
Xfd._6515_ fd._1692_ fd._1491_ VGND VGND VPWR VPWR fd._1694_ sky130_fd_sc_hd__nand2_1
XFILLER_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7495_ fd._2735_ VGND VGND VPWR VPWR fd._2772_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_114_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6446_ fd._1613_ fd._1614_ fd._1617_ VGND VGND VPWR VPWR fd._1618_ sky130_fd_sc_hd__mux2_2
XFILLER_25_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_283_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6377_ fd._0662_ fd._1540_ VGND VGND VPWR VPWR fd._1542_ sky130_fd_sc_hd__nand2_1
XFILLER_151_1489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8116_ fd._3431_ VGND VGND VPWR VPWR fd.ec\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_186_1519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5328_ fd._0000_ fd._0196_ fd._0198_ VGND VGND VPWR VPWR fd._0388_ sky130_fd_sc_hd__a21o_1
XFILLER_243_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8047_ fd._3378_ fd._3241_ VGND VGND VPWR VPWR fd._3379_ sky130_fd_sc_hd__nor2_1
XFILLER_252_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5259_ fd._3883_ VGND VGND VPWR VPWR fd._0312_ sky130_fd_sc_hd__inv_2
XFILLER_24_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_1503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_8428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_258_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_273_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_267_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_259_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput17 io_in[24] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput28 io_in[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_4
XFILLER_239_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4630_ fd.b\[11\] fd._3553_ fd._3554_ VGND VGND VPWR VPWR fd._3724_ sky130_fd_sc_hd__nand3_1
XFILLER_237_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_8962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_8984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._4561_ fd._3654_ VGND VGND VPWR VPWR fd._3655_ sky130_fd_sc_hd__inv_2
XFILLER_174_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_269_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6300_ fd._1416_ fd._1359_ fd._1415_ VGND VGND VPWR VPWR fd._1457_ sky130_fd_sc_hd__o21bai_1
XFILLER_46_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7280_ fd._2374_ fd._2383_ VGND VGND VPWR VPWR fd._2535_ sky130_fd_sc_hd__nand2_1
Xfd._4492_ fd._3585_ fd._2980_ VGND VGND VPWR VPWR fd._3586_ sky130_fd_sc_hd__xor2_1
XFILLER_113_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6231_ fd._1378_ fd._1380_ VGND VGND VPWR VPWR fd._1381_ sky130_fd_sc_hd__xnor2_1
XFILLER_77_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6162_ fd._1156_ fd._1160_ VGND VGND VPWR VPWR fd._1305_ sky130_fd_sc_hd__xor2_1
XFILLER_4_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5113_ fd._0150_ fd._4025_ VGND VGND VPWR VPWR fd._0151_ sky130_fd_sc_hd__xnor2_1
XFILLER_4_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6093_ fd._1146_ VGND VGND VPWR VPWR fd._1229_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_185_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5044_ fd._0074_ VGND VGND VPWR VPWR fd._0075_ sky130_fd_sc_hd__inv_2
XFILLER_209_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_1495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6995_ fd._2212_ fd._2213_ fd._2219_ fd._2220_ VGND VGND VPWR VPWR fd._2222_ sky130_fd_sc_hd__a31o_1
XFILLER_146_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_1700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5946_ fd._1063_ fd._1067_ fd._1047_ VGND VGND VPWR VPWR fd._1068_ sky130_fd_sc_hd__mux2_1
XFILLER_174_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5877_ fd._0837_ VGND VGND VPWR VPWR fd._0992_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_157_1610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7616_ fd._2900_ fd._2904_ fd._2875_ VGND VGND VPWR VPWR fd._2905_ sky130_fd_sc_hd__mux2_1
Xfd._4828_ fd._3832_ fd._3920_ fd._3921_ VGND VGND VPWR VPWR fd._3922_ sky130_fd_sc_hd__a21oi_1
XFILLER_270_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_249_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7547_ fd._2465_ fd._2828_ VGND VGND VPWR VPWR fd._2829_ sky130_fd_sc_hd__or2_1
XFILLER_130_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4759_ fd._3847_ fd._3851_ fd._3852_ VGND VGND VPWR VPWR fd._3853_ sky130_fd_sc_hd__a21o_1
XFILLER_170_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_275_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7478_ fd._1764_ fd._2623_ VGND VGND VPWR VPWR fd._2753_ sky130_fd_sc_hd__nor2_1
XFILLER_151_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6429_ fd._1558_ fd._1566_ fd._1596_ fd._1598_ fd._1555_ VGND VGND VPWR VPWR fd._1599_
+ sky130_fd_sc_hd__a311o_1
XFILLER_29_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_272_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_260_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_251_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_1671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_247_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_275_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_263_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5800_ fd._0904_ fd._0906_ VGND VGND VPWR VPWR fd._0907_ sky130_fd_sc_hd__xnor2_1
XFILLER_141_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_227_ fd.c\[19\] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_1
XFILLER_156_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6780_ fd._1956_ fd._1966_ fd._1982_ fd._1983_ fd._1984_ VGND VGND VPWR VPWR fd._1985_
+ sky130_fd_sc_hd__o311a_1
XFILLER_128_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5731_ fd._0638_ fd._0830_ VGND VGND VPWR VPWR fd._0831_ sky130_fd_sc_hd__nand2_1
XFILLER_183_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_256_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._5662_ fd._0653_ fd._0749_ fd._0754_ VGND VGND VPWR VPWR fd._0755_ sky130_fd_sc_hd__a21o_2
XTAP_8770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7401_ fd._2738_ fd._2667_ VGND VGND VPWR VPWR fd._2668_ sky130_fd_sc_hd__xnor2_1
XFILLER_98_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4613_ fd._3663_ fd._3706_ VGND VGND VPWR VPWR fd._3707_ sky130_fd_sc_hd__nand2_1
XFILLER_217_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5593_ fd._0677_ fd._0678_ VGND VGND VPWR VPWR fd._0679_ sky130_fd_sc_hd__xnor2_1
XFILLER_152_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_285_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7332_ fd._1797_ fd._2590_ VGND VGND VPWR VPWR fd._2592_ sky130_fd_sc_hd__or2_1
XFILLER_112_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4544_ fd._3555_ fd._3558_ VGND VGND VPWR VPWR fd._3638_ sky130_fd_sc_hd__nand2_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7263_ fd._1722_ fd._2514_ VGND VGND VPWR VPWR fd._2516_ sky130_fd_sc_hd__and2_1
XFILLER_117_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4475_ fd._0967_ fd._3568_ VGND VGND VPWR VPWR fd._3569_ sky130_fd_sc_hd__xnor2_1
XFILLER_78_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_250_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6214_ fd._1188_ VGND VGND VPWR VPWR fd._1362_ sky130_fd_sc_hd__clkinv_2
XFILLER_93_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7194_ fd._2223_ fd._2227_ VGND VGND VPWR VPWR fd._2440_ sky130_fd_sc_hd__nand2_1
XFILLER_265_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6145_ fd._1223_ fd._1285_ VGND VGND VPWR VPWR fd._1287_ sky130_fd_sc_hd__nor2_1
XFILLER_267_1660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_281_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_267_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6076_ fd._3537_ VGND VGND VPWR VPWR fd._1211_ sky130_fd_sc_hd__buf_6
XFILLER_181_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5027_ fd._0016_ fd._0023_ fd._0056_ fd._0051_ fd._0024_ VGND VGND VPWR VPWR fd._0057_
+ sky130_fd_sc_hd__a2111o_1
XFILLER_90_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6978_ fd._2201_ fd._2202_ VGND VGND VPWR VPWR fd._2203_ sky130_fd_sc_hd__nor2_1
XFILLER_159_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_1530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5929_ fd._0860_ VGND VGND VPWR VPWR fd._1049_ sky130_fd_sc_hd__clkinv_2
XFILLER_107_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_270_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_1659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_276_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_271_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_245_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_281_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_1398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_1406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_1439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_8066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4260_ fd._0219_ fd._1825_ VGND VGND VPWR VPWR fd._2045_ sky130_fd_sc_hd__nor2_1
XFILLER_207_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4191_ fd._1275_ VGND VGND VPWR VPWR fd._1286_ sky130_fd_sc_hd__buf_6
XFILLER_263_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7950_ fd._3169_ fd._3271_ VGND VGND VPWR VPWR fd._3272_ sky130_fd_sc_hd__nand2_1
XFILLER_91_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6901_ fd._2011_ fd._2010_ VGND VGND VPWR VPWR fd._2118_ sky130_fd_sc_hd__and2b_1
Xfd._7881_ fd._2326_ fd._3194_ VGND VGND VPWR VPWR fd._3196_ sky130_fd_sc_hd__nor2_1
XFILLER_31_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_1552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6832_ fd._1632_ fd._2041_ VGND VGND VPWR VPWR fd._2042_ sky130_fd_sc_hd__nand2_1
XFILLER_89_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6763_ fd._1958_ fd._1965_ VGND VGND VPWR VPWR fd._1966_ sky130_fd_sc_hd__and2_1
XFILLER_7_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_258_1659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5714_ fd._0262_ fd._0629_ VGND VGND VPWR VPWR fd._0812_ sky130_fd_sc_hd__or2_1
XFILLER_144_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6694_ fd._1889_ VGND VGND VPWR VPWR fd._1890_ sky130_fd_sc_hd__clkinvlp_2
XTAP_9290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_256_1383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5645_ fd._1308_ fd._0735_ VGND VGND VPWR VPWR fd._0737_ sky130_fd_sc_hd__or2_1
XFILLER_131_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_258_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5576_ fd._3833_ fd._0660_ VGND VGND VPWR VPWR fd._0661_ sky130_fd_sc_hd__or2_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_1670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7315_ fd._2571_ fd._2572_ VGND VGND VPWR VPWR fd._2574_ sky130_fd_sc_hd__nor2_1
XFILLER_112_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4527_ fd._3156_ fd._3178_ VGND VGND VPWR VPWR fd._3621_ sky130_fd_sc_hd__and2_1
XFILLER_230_1523 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_285_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7246_ fd._2426_ fd._2467_ fd._2480_ fd._2497_ VGND VGND VPWR VPWR fd._2498_ sky130_fd_sc_hd__or4_4
XFILLER_2_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4458_ fd._2243_ fd._3551_ fd._3211_ VGND VGND VPWR VPWR fd._3552_ sky130_fd_sc_hd__mux2_1
XFILLER_39_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_281_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7177_ fd._2258_ fd._2421_ VGND VGND VPWR VPWR fd._2422_ sky130_fd_sc_hd__xor2_1
Xfd._4389_ fd.b\[13\] fd._3365_ VGND VGND VPWR VPWR fd._3439_ sky130_fd_sc_hd__and2_1
XFILLER_226_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6128_ fd._1090_ fd._1096_ VGND VGND VPWR VPWR fd._1268_ sky130_fd_sc_hd__or2_1
XFILLER_228_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._6059_ fd._1015_ fd._1019_ VGND VGND VPWR VPWR fd._1192_ sky130_fd_sc_hd__or2_1
XFILLER_250_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_263_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_266_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_274_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_276_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_277_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_257_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_1632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5430_ fd._0497_ fd._0499_ fd._0425_ VGND VGND VPWR VPWR fd._0500_ sky130_fd_sc_hd__mux2_1
XTAP_7173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5361_ fd._0280_ fd._0416_ fd._0420_ fd._0423_ VGND VGND VPWR VPWR fd._0424_ sky130_fd_sc_hd__a31o_1
XTAP_6483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_269_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_255_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7100_ fd._2328_ fd._2336_ VGND VGND VPWR VPWR fd._2337_ sky130_fd_sc_hd__or2_1
XFILLER_83_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4312_ fd._0681_ fd._2606_ VGND VGND VPWR VPWR fd._2617_ sky130_fd_sc_hd__xnor2_1
XFILLER_212_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._8080_ fd._2020_ fd._2238_ fd._3398_ VGND VGND VPWR VPWR fd._3407_ sky130_fd_sc_hd__mux2_1
XFILLER_62_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5292_ fd._0343_ fd._0347_ VGND VGND VPWR VPWR fd._0348_ sky130_fd_sc_hd__nand2_1
XTAP_5793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._7031_ fd._1286_ fd._2260_ VGND VGND VPWR VPWR fd._2261_ sky130_fd_sc_hd__nand2_1
XFILLER_85_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4243_ fd.a\[2\] VGND VGND VPWR VPWR fd._1858_ sky130_fd_sc_hd__clkinv_2
XFILLER_209_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4174_ fd._1088_ fd.a\[20\] VGND VGND VPWR VPWR fd._1099_ sky130_fd_sc_hd__nor2_1
XFILLER_250_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_250_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7933_ fd._2863_ fd._3252_ VGND VGND VPWR VPWR fd._3253_ sky130_fd_sc_hd__or2_1
XFILLER_203_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7864_ fd._2142_ fd._3158_ fd._3175_ fd._3176_ VGND VGND VPWR VPWR fd._3177_ sky130_fd_sc_hd__a211oi_2
XFILLER_121_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_258_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6815_ fd._2017_ fd._1912_ VGND VGND VPWR VPWR fd._2024_ sky130_fd_sc_hd__xor2_1
XFILLER_145_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_258_1434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7795_ fd._2896_ fd._3100_ VGND VGND VPWR VPWR fd._3102_ sky130_fd_sc_hd__xnor2_1
XFILLER_8_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6746_ fd._1947_ VGND VGND VPWR VPWR fd._1948_ sky130_fd_sc_hd__inv_2
XFILLER_145_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_271_1612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6677_ fd._0716_ VGND VGND VPWR VPWR fd._1872_ sky130_fd_sc_hd__buf_6
XFILLER_154_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_1530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5628_ fd._0717_ fd._0661_ VGND VGND VPWR VPWR fd._0718_ sky130_fd_sc_hd__nand2_1
XFILLER_119_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_258_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_285_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5559_ fd._0427_ fd._0622_ VGND VGND VPWR VPWR fd._0642_ sky130_fd_sc_hd__nor2_1
XFILLER_140_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7229_ fd._2476_ fd._2478_ VGND VGND VPWR VPWR fd._2479_ sky130_fd_sc_hd__and2_1
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_281_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_276_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_269_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4930_ fd._3708_ fd._4023_ VGND VGND VPWR VPWR fd._4024_ sky130_fd_sc_hd__or2_1
XFILLER_125_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._4861_ fd._3781_ fd._3944_ fd._3767_ VGND VGND VPWR VPWR fd._3955_ sky130_fd_sc_hd__a21o_1
XFILLER_195_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6600_ fd._1784_ fd._1729_ fd._1783_ VGND VGND VPWR VPWR fd._1787_ sky130_fd_sc_hd__o21bai_1
XFILLER_86_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7580_ fd._2862_ fd._2864_ VGND VGND VPWR VPWR fd._2865_ sky130_fd_sc_hd__nor2_1
XFILLER_127_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4792_ fd._3669_ fd._3857_ VGND VGND VPWR VPWR fd._3886_ sky130_fd_sc_hd__or2_1
XFILLER_142_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_275_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6531_ fd._1643_ fd._1631_ VGND VGND VPWR VPWR fd._1711_ sky130_fd_sc_hd__and2b_1
XFILLER_153_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6462_ fd._1633_ fd._1634_ fd._1617_ VGND VGND VPWR VPWR fd._1635_ sky130_fd_sc_hd__or3b_1
XFILLER_214_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8201_ net66 fd.ec\[2\] VGND VGND VPWR VPWR fd.c\[25\] sky130_fd_sc_hd__dfxtp_1
Xfd._5413_ fd._0469_ fd._0476_ fd._0478_ fd._0480_ fd._0454_ VGND VGND VPWR VPWR fd._0481_
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_136_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6393_ fd._0807_ VGND VGND VPWR VPWR fd._1559_ sky130_fd_sc_hd__buf_6
XFILLER_256_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8132_ fd._3436_ fd._3446_ VGND VGND VPWR VPWR fd._3447_ sky130_fd_sc_hd__nand2_1
Xfd._5344_ fd._0404_ fd._0210_ VGND VGND VPWR VPWR fd._0405_ sky130_fd_sc_hd__nor2_1
XFILLER_23_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_282_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8063_ fd._1231_ fd._3395_ VGND VGND VPWR VPWR fd._3396_ sky130_fd_sc_hd__and2_1
Xfd._5275_ fd._0311_ fd._0317_ fd._0328_ fd._0309_ VGND VGND VPWR VPWR fd._0330_ sky130_fd_sc_hd__o31a_1
XFILLER_282_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7014_ fd._2036_ fd._2238_ VGND VGND VPWR VPWR fd._2242_ sky130_fd_sc_hd__nor2_1
XFILLER_63_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4226_ fd._0461_ fd._1660_ VGND VGND VPWR VPWR fd._1671_ sky130_fd_sc_hd__nand2_1
XFILLER_184_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_263_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_282_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_251_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4157_ fd._0846_ fd.a\[11\] fd._0890_ fd._0901_ VGND VGND VPWR VPWR fd._0912_
+ sky130_fd_sc_hd__o22ai_1
XFILLER_211_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4088_ fd._0076_ fd.a\[18\] VGND VGND VPWR VPWR fd._0153_ sky130_fd_sc_hd__nand2_1
XFILLER_143_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7916_ fd._3231_ fd._3234_ fd._3077_ VGND VGND VPWR VPWR fd._3235_ sky130_fd_sc_hd__mux2_1
XFILLER_143_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7847_ fd._2763_ fd._2956_ VGND VGND VPWR VPWR fd._3159_ sky130_fd_sc_hd__nor2_1
XFILLER_192_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7778_ fd._2893_ fd._3016_ VGND VGND VPWR VPWR fd._3083_ sky130_fd_sc_hd__or2b_1
XFILLER_145_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6729_ fd._1927_ fd._1928_ VGND VGND VPWR VPWR fd._1929_ sky130_fd_sc_hd__xnor2_1
XFILLER_195_1598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_259_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_265_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_276_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_269_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5060_ fd._4017_ fd._0092_ VGND VGND VPWR VPWR fd._0093_ sky130_fd_sc_hd__nand2_1
XTAP_3473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_283_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5962_ fd._0919_ fd._1084_ VGND VGND VPWR VPWR fd._1085_ sky130_fd_sc_hd__xnor2_1
XFILLER_158_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7701_ fd._1645_ fd._2992_ fd._2997_ VGND VGND VPWR VPWR fd._2998_ sky130_fd_sc_hd__mux2_1
XFILLER_31_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4913_ fd.b\[1\] fd._3875_ VGND VGND VPWR VPWR fd._4007_ sky130_fd_sc_hd__and2_1
Xfd._5893_ fd._0826_ VGND VGND VPWR VPWR fd._1009_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_173_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4844_ fd._3937_ VGND VGND VPWR VPWR fd._3938_ sky130_fd_sc_hd__inv_2
Xfd._7632_ fd._2533_ fd._2741_ VGND VGND VPWR VPWR fd._2922_ sky130_fd_sc_hd__or2_1
XFILLER_127_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_project_wrapper_120 VGND VGND VPWR VPWR user_project_wrapper_120/HI io_out[36]
+ sky130_fd_sc_hd__conb_1
XFILLER_259_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_255_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_project_wrapper_131 VGND VGND VPWR VPWR user_project_wrapper_131/HI la_data_out[9]
+ sky130_fd_sc_hd__conb_1
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_project_wrapper_142 VGND VGND VPWR VPWR user_project_wrapper_142/HI la_data_out[20]
+ sky130_fd_sc_hd__conb_1
XFILLER_99_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_153 VGND VGND VPWR VPWR user_project_wrapper_153/HI la_data_out[31]
+ sky130_fd_sc_hd__conb_1
Xfd._4775_ fd.b\[3\] VGND VGND VPWR VPWR fd._3869_ sky130_fd_sc_hd__buf_6
XFILLER_217_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7563_ fd._2844_ fd._2845_ VGND VGND VPWR VPWR fd._2846_ sky130_fd_sc_hd__and2b_1
Xuser_project_wrapper_164 VGND VGND VPWR VPWR user_project_wrapper_164/HI la_data_out[42]
+ sky130_fd_sc_hd__conb_1
XFILLER_142_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_project_wrapper_175 VGND VGND VPWR VPWR user_project_wrapper_175/HI la_data_out[53]
+ sky130_fd_sc_hd__conb_1
XFILLER_114_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_186 VGND VGND VPWR VPWR user_project_wrapper_186/HI la_data_out[64]
+ sky130_fd_sc_hd__conb_1
XFILLER_64_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6514_ fd._1482_ fd._1488_ fd._1492_ VGND VGND VPWR VPWR fd._1692_ sky130_fd_sc_hd__a21o_1
XFILLER_130_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_project_wrapper_197 VGND VGND VPWR VPWR user_project_wrapper_197/HI la_data_out[75]
+ sky130_fd_sc_hd__conb_1
XFILLER_269_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7494_ fd._0312_ fd._2743_ fd._2750_ fd._2768_ fd._2769_ VGND VGND VPWR VPWR fd._2770_
+ sky130_fd_sc_hd__a221o_1
XFILLER_64_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6445_ fd._1615_ VGND VGND VPWR VPWR fd._1617_ sky130_fd_sc_hd__buf_6
XFILLER_68_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_256_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._6376_ fd._0662_ fd._1540_ VGND VGND VPWR VPWR fd._1541_ sky130_fd_sc_hd__or2_1
XFILLER_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8115_ fd._3428_ fd._3429_ VGND VGND VPWR VPWR fd._3431_ sky130_fd_sc_hd__or2_1
Xfd._5327_ fd._0288_ fd._0386_ fd._0282_ fd._1264_ VGND VGND VPWR VPWR fd._0387_ sky130_fd_sc_hd__a22o_1
XFILLER_266_1511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8046_ fd._3095_ VGND VGND VPWR VPWR fd._3378_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_224_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5258_ fd._0309_ fd._0310_ VGND VGND VPWR VPWR fd._0311_ sky130_fd_sc_hd__nand2_1
XFILLER_3_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4209_ fd._1462_ fd._1473_ fd._0527_ VGND VGND VPWR VPWR fd._1484_ sky130_fd_sc_hd__o21ai_1
XFILLER_262_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5189_ fd._0228_ fd._0234_ fd._0233_ VGND VGND VPWR VPWR fd._0235_ sky130_fd_sc_hd__a21o_1
XFILLER_212_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1662 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_277_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_258_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_262_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_284_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput18 io_in[25] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput29 io_in[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_4
XFILLER_182_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4560_ fd._3469_ fd._3653_ VGND VGND VPWR VPWR fd._3654_ sky130_fd_sc_hd__nor2_1
XFILLER_233_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4491_ fd._2705_ fd._2672_ fd._2694_ VGND VGND VPWR VPWR fd._3585_ sky130_fd_sc_hd__a21oi_1
XFILLER_133_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6230_ fd._1205_ fd._1379_ VGND VGND VPWR VPWR fd._1380_ sky130_fd_sc_hd__nand2_1
XFILLER_120_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_280_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6161_ fd._0482_ VGND VGND VPWR VPWR fd._1304_ sky130_fd_sc_hd__buf_6
XFILLER_225_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5112_ fd._3980_ fd._3979_ fd._0149_ VGND VGND VPWR VPWR fd._0150_ sky130_fd_sc_hd__o21a_1
XFILLER_93_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_280_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_283_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6092_ fd._1177_ fd._1227_ VGND VGND VPWR VPWR fd._1228_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5043_ fd._1253_ fd._0073_ VGND VGND VPWR VPWR fd._0074_ sky130_fd_sc_hd__or2_1
XFILLER_59_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_244_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6994_ fd._1656_ fd._2218_ VGND VGND VPWR VPWR fd._2220_ sky130_fd_sc_hd__nor2_1
XFILLER_14_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5945_ fd._1065_ fd._0977_ VGND VGND VPWR VPWR fd._1067_ sky130_fd_sc_hd__xnor2_1
XFILLER_158_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5876_ fd._0819_ fd._0836_ fd._0817_ VGND VGND VPWR VPWR fd._0991_ sky130_fd_sc_hd__a21o_1
XFILLER_174_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_259_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._7615_ fd._2902_ fd._2779_ VGND VGND VPWR VPWR fd._2904_ sky130_fd_sc_hd__xnor2_1
Xfd._4827_ fd._3646_ fd._3827_ VGND VGND VPWR VPWR fd._3921_ sky130_fd_sc_hd__and2_1
XFILLER_161_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4758_ fd._3469_ fd._3845_ VGND VGND VPWR VPWR fd._3852_ sky130_fd_sc_hd__and2_1
XFILLER_216_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7546_ fd._2644_ fd._2827_ fd._2813_ VGND VGND VPWR VPWR fd._2828_ sky130_fd_sc_hd__mux2_1
XFILLER_114_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_275_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_257_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4689_ fd._3777_ fd._3779_ fd._3782_ VGND VGND VPWR VPWR fd._3783_ sky130_fd_sc_hd__or3_1
Xfd._7477_ fd._2556_ fd._2670_ fd._2675_ VGND VGND VPWR VPWR fd._2752_ sky130_fd_sc_hd__nand3_1
XFILLER_130_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6428_ fd._1219_ fd._1597_ VGND VGND VPWR VPWR fd._1598_ sky130_fd_sc_hd__nor2_1
XFILLER_112_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_283_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6359_ fd._0786_ fd._1521_ VGND VGND VPWR VPWR fd._1522_ sky130_fd_sc_hd__or2_1
XFILLER_95_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_272_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8029_ fd._3331_ fd._3330_ fd._3322_ fd._3358_ VGND VGND VPWR VPWR fd._3359_ sky130_fd_sc_hd__o31a_1
XFILLER_24_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_273_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_277_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_219_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_262_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_226_ fd.c\[18\] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_1
XFILLER_54_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5730_ fd._0828_ fd._0801_ fd._0672_ fd._0829_ VGND VGND VPWR VPWR fd._0830_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_7_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5661_ fd._0594_ fd._0753_ VGND VGND VPWR VPWR fd._0754_ sky130_fd_sc_hd__xnor2_1
XFILLER_143_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4612_ fd._2155_ fd._3661_ VGND VGND VPWR VPWR fd._3706_ sky130_fd_sc_hd__nand2_1
XFILLER_252_1407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7400_ fd._2493_ fd._2666_ fd._2623_ VGND VGND VPWR VPWR fd._2667_ sky130_fd_sc_hd__mux2_2
XTAP_8782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5592_ fd._0520_ fd._0522_ VGND VGND VPWR VPWR fd._0678_ sky130_fd_sc_hd__or2_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4543_ fd._1253_ fd._3636_ VGND VGND VPWR VPWR fd._3637_ sky130_fd_sc_hd__or2_1
XFILLER_170_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7331_ fd._1797_ fd._2590_ VGND VGND VPWR VPWR fd._2591_ sky130_fd_sc_hd__nand2_1
XFILLER_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_257_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7262_ fd._1722_ fd._2514_ VGND VGND VPWR VPWR fd._2515_ sky130_fd_sc_hd__nor2_1
Xfd._4474_ fd._2529_ fd._3567_ fd._3222_ VGND VGND VPWR VPWR fd._3568_ sky130_fd_sc_hd__mux2_1
XFILLER_239_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_272_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6213_ fd._1359_ fd._1360_ VGND VGND VPWR VPWR fd._1361_ sky130_fd_sc_hd__nor2_1
XFILLER_281_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7193_ fd._1685_ fd._2438_ VGND VGND VPWR VPWR fd._2439_ sky130_fd_sc_hd__or2_1
XFILLER_113_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6144_ fd._4055_ fd._1131_ VGND VGND VPWR VPWR fd._1285_ sky130_fd_sc_hd__xnor2_1
XFILLER_4_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_225_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6075_ fd._0985_ fd._1206_ fd._1208_ VGND VGND VPWR VPWR fd._1210_ sky130_fd_sc_hd__o21bai_2
XFILLER_234_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5026_ fd._0035_ fd._0055_ VGND VGND VPWR VPWR fd._0056_ sky130_fd_sc_hd__nand2_1
XFILLER_181_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6977_ fd._1600_ fd._2200_ VGND VGND VPWR VPWR fd._2202_ sky130_fd_sc_hd__nor2_1
XFILLER_200_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5928_ fd._0855_ fd._1045_ fd._1047_ VGND VGND VPWR VPWR fd._1048_ sky130_fd_sc_hd__mux2_1
XFILLER_190_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_274_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5859_ fd._0743_ fd._0971_ fd._0849_ VGND VGND VPWR VPWR fd._0972_ sky130_fd_sc_hd__mux2_1
XFILLER_200_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7529_ fd._1685_ fd._2808_ VGND VGND VPWR VPWR fd._2809_ sky130_fd_sc_hd__nor2_1
XTAP_5419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_268_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_268_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_260_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_262_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_8089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_273_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4190_ fd._1264_ VGND VGND VPWR VPWR fd._1275_ sky130_fd_sc_hd__buf_6
XFILLER_5_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6900_ fd._1918_ fd._2015_ fd._2116_ VGND VGND VPWR VPWR fd._2117_ sky130_fd_sc_hd__mux2_1
XFILLER_148_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7880_ fd._2326_ fd._3194_ VGND VGND VPWR VPWR fd._3195_ sky130_fd_sc_hd__nand2_1
XFILLER_19_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6831_ fd._1906_ fd._2040_ fd._2020_ VGND VGND VPWR VPWR fd._2041_ sky130_fd_sc_hd__mux2_2
XFILLER_15_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_209_ fd.c\[1\] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_1
XFILLER_15_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6762_ fd._1959_ fd._1964_ fd._1916_ VGND VGND VPWR VPWR fd._1965_ sky130_fd_sc_hd__mux2_1
XFILLER_128_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5713_ fd._0638_ fd._0636_ fd._0639_ VGND VGND VPWR VPWR fd._0811_ sky130_fd_sc_hd__o21ai_1
XFILLER_183_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._6693_ fd._1864_ fd._1888_ VGND VGND VPWR VPWR fd._1889_ sky130_fd_sc_hd__nor2_1
XFILLER_144_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_256_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._5644_ fd._0732_ fd._0733_ fd._0672_ fd._0734_ VGND VGND VPWR VPWR fd._0735_ sky130_fd_sc_hd__o31a_1
XFILLER_154_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5575_ fd._0546_ fd._0658_ fd._0614_ VGND VGND VPWR VPWR fd._0660_ sky130_fd_sc_hd__mux2_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7314_ fd._2566_ fd._2570_ VGND VGND VPWR VPWR fd._2572_ sky130_fd_sc_hd__nor2_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4526_ fd._3189_ fd._3156_ fd._3178_ VGND VGND VPWR VPWR fd._3620_ sky130_fd_sc_hd__a21oi_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_226_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4457_ fd._2298_ fd._3550_ VGND VGND VPWR VPWR fd._3551_ sky130_fd_sc_hd__xnor2_1
XFILLER_187_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._7245_ fd._2489_ fd._2495_ VGND VGND VPWR VPWR fd._2497_ sky130_fd_sc_hd__nand2_1
XFILLER_38_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1579 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4388_ fd.b\[15\] fd._3277_ VGND VGND VPWR VPWR fd._3430_ sky130_fd_sc_hd__xnor2_1
XFILLER_199_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7176_ fd._2261_ fd._2290_ VGND VGND VPWR VPWR fd._2421_ sky130_fd_sc_hd__nand2_1
XFILLER_113_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_281_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_263_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6127_ fd._1258_ fd._1263_ fd._1266_ fd._1256_ VGND VGND VPWR VPWR fd._1267_ sky130_fd_sc_hd__o31a_1
XFILLER_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6058_ fd._1025_ fd._1028_ VGND VGND VPWR VPWR fd._1191_ sky130_fd_sc_hd__nand2_1
XFILLER_62_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5009_ fd._3773_ fd._3966_ VGND VGND VPWR VPWR fd._0037_ sky130_fd_sc_hd__or2_1
XFILLER_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_1503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_270_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_282_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_268_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5360_ fd._0271_ fd._0277_ fd._0422_ VGND VGND VPWR VPWR fd._0423_ sky130_fd_sc_hd__o21ai_1
XFILLER_27_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_251_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4311_ fd._0703_ fd._2518_ fd._0692_ VGND VGND VPWR VPWR fd._2606_ sky130_fd_sc_hd__a21o_1
XFILLER_255_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5291_ fd._0344_ fd._0346_ fd._0269_ VGND VGND VPWR VPWR fd._0347_ sky130_fd_sc_hd__mux2_1
XTAP_5783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4242_ fd._1836_ VGND VGND VPWR VPWR fd._1847_ sky130_fd_sc_hd__inv_2
XFILLER_224_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7030_ fd._2072_ fd._2259_ fd._2238_ VGND VGND VPWR VPWR fd._2260_ sky130_fd_sc_hd__mux2_1
XFILLER_91_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_263_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4173_ fd.b\[20\] VGND VGND VPWR VPWR fd._1088_ sky130_fd_sc_hd__inv_2
XFILLER_211_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_260_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7932_ fd._3226_ fd._3251_ fd._3240_ VGND VGND VPWR VPWR fd._3252_ sky130_fd_sc_hd__mux2_1
XFILLER_31_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7863_ fd._2533_ fd._3151_ VGND VGND VPWR VPWR fd._3176_ sky130_fd_sc_hd__nor2_1
XFILLER_31_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6814_ fd._1823_ VGND VGND VPWR VPWR fd._2022_ sky130_fd_sc_hd__clkinv_2
XFILLER_157_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7794_ fd._2990_ fd._2989_ fd._3076_ VGND VGND VPWR VPWR fd._3100_ sky130_fd_sc_hd__nand3b_1
XFILLER_145_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_258_1446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._6745_ fd._1755_ fd._1945_ fd._1916_ VGND VGND VPWR VPWR fd._1947_ sky130_fd_sc_hd__mux2_1
XFILLER_156_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6676_ fd._1870_ VGND VGND VPWR VPWR fd._1871_ sky130_fd_sc_hd__clkinv_4
XFILLER_98_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_258_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5627_ fd._0716_ fd._0660_ VGND VGND VPWR VPWR fd._0717_ sky130_fd_sc_hd__nand2_1
XFILLER_154_1444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_258_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_274_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5558_ fd._0630_ fd._0640_ VGND VGND VPWR VPWR fd._0641_ sky130_fd_sc_hd__and2_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4509_ fd._2870_ fd._3602_ fd._3222_ VGND VGND VPWR VPWR fd._3603_ sky130_fd_sc_hd__mux2_1
XFILLER_227_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_285_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5489_ fd._0292_ fd._0361_ fd._0368_ VGND VGND VPWR VPWR fd._0565_ sky130_fd_sc_hd__and3_1
XFILLER_22_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7228_ fd._2477_ VGND VGND VPWR VPWR fd._2478_ sky130_fd_sc_hd__inv_2
XFILLER_2_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_282_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7159_ fd._2211_ fd._2401_ fd._2323_ VGND VGND VPWR VPWR fd._2402_ sky130_fd_sc_hd__mux2_1
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_1588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4860_ fd._3937_ fd._3942_ fd._3953_ VGND VGND VPWR VPWR fd._3954_ sky130_fd_sc_hd__a21o_2
XFILLER_200_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4791_ fd._3868_ fd._3874_ fd._3881_ fd._3882_ fd._3884_ VGND VGND VPWR VPWR fd._3885_
+ sky130_fd_sc_hd__a311o_1
XFILLER_181_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6530_ fd._1632_ fd._1636_ VGND VGND VPWR VPWR fd._1710_ sky130_fd_sc_hd__or2_1
XFILLER_142_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_1452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_253_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6461_ fd._1434_ fd._1500_ fd._1502_ VGND VGND VPWR VPWR fd._1634_ sky130_fd_sc_hd__and3_1
XFILLER_171_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._8200_ net66 fd.ec\[1\] VGND VGND VPWR VPWR fd.c\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_256_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5412_ fd._0479_ fd._0468_ VGND VGND VPWR VPWR fd._0480_ sky130_fd_sc_hd__nand2_1
XFILLER_150_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._6392_ fd._1557_ VGND VGND VPWR VPWR fd._1558_ sky130_fd_sc_hd__inv_2
XFILLER_171_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8131_ fd._3444_ fd._3445_ VGND VGND VPWR VPWR fd._3446_ sky130_fd_sc_hd__or2_1
XFILLER_231_1652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5343_ fd._0070_ VGND VGND VPWR VPWR fd._0404_ sky130_fd_sc_hd__inv_2
XFILLER_209_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_255_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5274_ fd._0324_ fd._0325_ fd._0326_ fd._0327_ VGND VGND VPWR VPWR fd._0328_ sky130_fd_sc_hd__o211a_1
XFILLER_209_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8062_ fd._3264_ fd._3384_ fd._3394_ VGND VGND VPWR VPWR fd._3395_ sky130_fd_sc_hd__a21o_1
XFILLER_270_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_282_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4225_ fd._0230_ fd._1649_ VGND VGND VPWR VPWR fd._1660_ sky130_fd_sc_hd__nand2_1
Xfd._7013_ fd._2235_ fd._2110_ VGND VGND VPWR VPWR fd._2241_ sky130_fd_sc_hd__or2_1
XFILLER_58_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_282_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4156_ fd._0846_ fd.a\[11\] fd._0571_ VGND VGND VPWR VPWR fd._0901_ sky130_fd_sc_hd__a21o_1
XFILLER_225_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4087_ fd._0131_ fd.a\[19\] VGND VGND VPWR VPWR fd._0142_ sky130_fd_sc_hd__nand2_1
XFILLER_52_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7915_ fd._3037_ fd._3232_ VGND VGND VPWR VPWR fd._3234_ sky130_fd_sc_hd__xnor2_1
XFILLER_137_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7846_ fd._3153_ fd._3157_ fd._3075_ VGND VGND VPWR VPWR fd._3158_ sky130_fd_sc_hd__mux2_2
XFILLER_118_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_247_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7777_ fd._3009_ fd._3015_ fd._3017_ VGND VGND VPWR VPWR fd._3082_ sky130_fd_sc_hd__o21a_1
Xfd._4989_ fd._3580_ fd._0013_ VGND VGND VPWR VPWR fd._0015_ sky130_fd_sc_hd__nor2_1
XFILLER_160_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6728_ fd._1736_ fd._1777_ VGND VGND VPWR VPWR fd._1928_ sky130_fd_sc_hd__or2b_1
XFILLER_145_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._6659_ fd._1494_ fd._1851_ VGND VGND VPWR VPWR fd._1852_ sky130_fd_sc_hd__nand2_1
XFILLER_132_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_271_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_259_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_214_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_1545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_269_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_1656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5961_ fd._0929_ fd._0925_ VGND VGND VPWR VPWR fd._1084_ sky130_fd_sc_hd__nor2_1
XFILLER_144_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7700_ fd._1645_ fd._2996_ VGND VGND VPWR VPWR fd._2997_ sky130_fd_sc_hd__xnor2_1
Xfd._4912_ fd._3695_ fd._3788_ fd._3954_ fd._3958_ VGND VGND VPWR VPWR fd._4006_ sky130_fd_sc_hd__o211a_1
XFILLER_174_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._5892_ fd._0831_ fd._0833_ VGND VGND VPWR VPWR fd._1008_ sky130_fd_sc_hd__nand2_1
Xfd._7631_ fd._2750_ fd._2768_ fd._2769_ VGND VGND VPWR VPWR fd._2921_ sky130_fd_sc_hd__a21o_1
XFILLER_127_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._4843_ fd._3773_ fd._3789_ VGND VGND VPWR VPWR fd._3937_ sky130_fd_sc_hd__or2_1
XFILLER_31_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_project_wrapper_110 VGND VGND VPWR VPWR user_project_wrapper_110/HI io_oeb[32]
+ sky130_fd_sc_hd__conb_1
XFILLER_142_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_121 VGND VGND VPWR VPWR user_project_wrapper_121/HI io_out[37]
+ sky130_fd_sc_hd__conb_1
XFILLER_259_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_project_wrapper_132 VGND VGND VPWR VPWR user_project_wrapper_132/HI la_data_out[10]
+ sky130_fd_sc_hd__conb_1
XFILLER_66_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7562_ fd._1242_ fd._2843_ VGND VGND VPWR VPWR fd._2845_ sky130_fd_sc_hd__nand2_1
Xuser_project_wrapper_143 VGND VGND VPWR VPWR user_project_wrapper_143/HI la_data_out[21]
+ sky130_fd_sc_hd__conb_1
Xfd._4774_ fd._0450_ fd._3867_ VGND VGND VPWR VPWR fd._3868_ sky130_fd_sc_hd__xnor2_1
Xuser_project_wrapper_154 VGND VGND VPWR VPWR user_project_wrapper_154/HI la_data_out[32]
+ sky130_fd_sc_hd__conb_1
XFILLER_47_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_165 VGND VGND VPWR VPWR user_project_wrapper_165/HI la_data_out[43]
+ sky130_fd_sc_hd__conb_1
XFILLER_217_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_project_wrapper_176 VGND VGND VPWR VPWR user_project_wrapper_176/HI la_data_out[54]
+ sky130_fd_sc_hd__conb_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6513_ fd._1443_ VGND VGND VPWR VPWR fd._1691_ sky130_fd_sc_hd__clkinv_2
Xuser_project_wrapper_187 VGND VGND VPWR VPWR user_project_wrapper_187/HI la_data_out[65]
+ sky130_fd_sc_hd__conb_1
Xfd._7493_ fd._2142_ fd._2748_ VGND VGND VPWR VPWR fd._2769_ sky130_fd_sc_hd__and2_1
XFILLER_114_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_project_wrapper_198 VGND VGND VPWR VPWR user_project_wrapper_198/HI la_data_out[76]
+ sky130_fd_sc_hd__conb_1
XFILLER_99_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6444_ fd._1533_ VGND VGND VPWR VPWR fd._1615_ sky130_fd_sc_hd__buf_6
XFILLER_64_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_256_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6375_ fd._1410_ fd._1538_ fd._1533_ VGND VGND VPWR VPWR fd._1540_ sky130_fd_sc_hd__mux2_1
XFILLER_256_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8114_ fd._1231_ fd._3427_ VGND VGND VPWR VPWR fd._3429_ sky130_fd_sc_hd__and2_1
XFILLER_3_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5326_ fd._0375_ fd._0379_ fd._0381_ fd._0385_ VGND VGND VPWR VPWR fd._0386_ sky130_fd_sc_hd__a211o_1
XFILLER_7_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_255_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_1523 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._8045_ fd._3206_ fd._3105_ fd._3122_ fd._3203_ VGND VGND VPWR VPWR fd._3377_ sky130_fd_sc_hd__nand4_1
Xfd._5257_ fd._3669_ fd._0308_ VGND VGND VPWR VPWR fd._0310_ sky130_fd_sc_hd__nand2_1
XFILLER_70_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4208_ fd._1385_ fd._0626_ fd._0604_ VGND VGND VPWR VPWR fd._1473_ sky130_fd_sc_hd__a21oi_1
XFILLER_24_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5188_ fd._0232_ fd._0233_ VGND VGND VPWR VPWR fd._0234_ sky130_fd_sc_hd__nor2_2
XFILLER_224_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_212_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4139_ fd._0692_ fd._0703_ VGND VGND VPWR VPWR fd._0714_ sky130_fd_sc_hd__and2b_1
XFILLER_211_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7829_ fd._2926_ fd._3138_ fd._3075_ VGND VGND VPWR VPWR fd._3139_ sky130_fd_sc_hd__mux2_1
XTAP_8419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_1330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_273_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_274_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_275_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_261_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_265_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_284_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_1632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput19 io_in[26] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_1
XFILLER_156_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_8953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_269_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4490_ fd._3578_ fd._3583_ VGND VGND VPWR VPWR fd._3584_ sky130_fd_sc_hd__xnor2_1
XFILLER_61_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_285_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6160_ fd._0207_ fd._1298_ fd._1302_ VGND VGND VPWR VPWR fd._1303_ sky130_fd_sc_hd__mux2_2
XFILLER_237_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_280_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5111_ fd._4027_ fd._0080_ VGND VGND VPWR VPWR fd._0149_ sky130_fd_sc_hd__or2_1
XFILLER_185_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6091_ fd._1218_ fd._1225_ fd._1226_ VGND VGND VPWR VPWR fd._1227_ sky130_fd_sc_hd__o21a_1
XFILLER_185_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5042_ fd._0072_ fd._0003_ fd._0067_ VGND VGND VPWR VPWR fd._0073_ sky130_fd_sc_hd__mux2_1
XTAP_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_283_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6993_ fd._1656_ fd._2218_ VGND VGND VPWR VPWR fd._2219_ sky130_fd_sc_hd__nand2_1
XFILLER_144_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5944_ fd._0974_ fd._1064_ fd._0884_ VGND VGND VPWR VPWR fd._1065_ sky130_fd_sc_hd__o21ba_1
XFILLER_179_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5875_ fd._0988_ VGND VGND VPWR VPWR fd._0990_ sky130_fd_sc_hd__clkinv_2
XFILLER_179_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_255_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7614_ fd._2785_ fd._2901_ fd._2725_ VGND VGND VPWR VPWR fd._2902_ sky130_fd_sc_hd__a21boi_1
Xfd._4826_ fd._3841_ fd._3916_ fd._3919_ fd._3839_ VGND VGND VPWR VPWR fd._3920_ sky130_fd_sc_hd__a211o_1
XFILLER_196_1683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_1634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_255_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7545_ fd._2823_ fd._2825_ VGND VGND VPWR VPWR fd._2827_ sky130_fd_sc_hd__xnor2_1
Xfd._4757_ fd._2155_ fd._3850_ VGND VGND VPWR VPWR fd._3851_ sky130_fd_sc_hd__or2_1
XFILLER_118_1629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7476_ fd._1958_ VGND VGND VPWR VPWR fd._2751_ sky130_fd_sc_hd__buf_6
Xfd._4688_ fd._3763_ fd._3781_ VGND VGND VPWR VPWR fd._3782_ sky130_fd_sc_hd__nand2_1
XFILLER_9_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_256_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6427_ fd._1546_ VGND VGND VPWR VPWR fd._1597_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_3_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_272_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6358_ fd._1333_ fd._1515_ fd._1423_ VGND VGND VPWR VPWR fd._1521_ sky130_fd_sc_hd__mux2_1
XFILLER_113_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5309_ fd._3917_ fd._0366_ VGND VGND VPWR VPWR fd._0367_ sky130_fd_sc_hd__nor2_1
XFILLER_260_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6289_ fd._1272_ VGND VGND VPWR VPWR fd._1445_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_266_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._8028_ fd._3318_ fd._3320_ VGND VGND VPWR VPWR fd._3358_ sky130_fd_sc_hd__nand2_1
XFILLER_64_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_262_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_1668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_8205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_277_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_259_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_270_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_262_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_243_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_225_ fd.c\[17\] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_1
XFILLER_15_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_1500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5660_ fd._0589_ fd._0752_ fd._0651_ VGND VGND VPWR VPWR fd._0753_ sky130_fd_sc_hd__mux2_1
XFILLER_48_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4611_ fd._0428_ fd._3704_ VGND VGND VPWR VPWR fd._3705_ sky130_fd_sc_hd__or2_1
XTAP_8772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_8783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._5591_ fd._0430_ fd._0447_ fd._0523_ VGND VGND VPWR VPWR fd._0677_ sky130_fd_sc_hd__a21o_1
XFILLER_139_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._7330_ fd._2587_ fd._2589_ fd._2506_ VGND VGND VPWR VPWR fd._2590_ sky130_fd_sc_hd__mux2_1
XFILLER_112_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4542_ fd._3568_ fd._3635_ fd._3625_ VGND VGND VPWR VPWR fd._3636_ sky130_fd_sc_hd__mux2_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7261_ fd._2512_ fd._2506_ fd._2513_ VGND VGND VPWR VPWR fd._2514_ sky130_fd_sc_hd__a21oi_1
XFILLER_117_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4473_ fd._2496_ fd._3566_ VGND VGND VPWR VPWR fd._3567_ sky130_fd_sc_hd__xnor2_1
XFILLER_66_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6212_ fd._1173_ fd._1357_ VGND VGND VPWR VPWR fd._1360_ sky130_fd_sc_hd__nor2_1
XFILLER_254_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._7192_ fd._2436_ fd._2323_ fd._2437_ VGND VGND VPWR VPWR fd._2438_ sky130_fd_sc_hd__a21oi_1
XFILLER_285_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_265_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_280_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6143_ fd._1127_ fd._1131_ VGND VGND VPWR VPWR fd._1284_ sky130_fd_sc_hd__xnor2_1
XFILLER_92_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_280_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6074_ fd._1059_ fd._1074_ fd._1167_ fd._1207_ fd._1200_ VGND VGND VPWR VPWR fd._1208_
+ sky130_fd_sc_hd__o311a_1
XTAP_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_263_1548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_1668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5025_ fd._0053_ fd._3967_ VGND VGND VPWR VPWR fd._0055_ sky130_fd_sc_hd__nor2_1
XFILLER_233_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6976_ fd._1600_ fd._2200_ VGND VGND VPWR VPWR fd._2201_ sky130_fd_sc_hd__and2_1
XFILLER_124_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5927_ fd._1046_ VGND VGND VPWR VPWR fd._1047_ sky130_fd_sc_hd__buf_6
XFILLER_174_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_274_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5858_ fd._0000_ fd._0744_ VGND VGND VPWR VPWR fd._0971_ sky130_fd_sc_hd__xnor2_1
XFILLER_161_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_255_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4809_ fd._3902_ fd._3653_ fd._3787_ VGND VGND VPWR VPWR fd._3903_ sky130_fd_sc_hd__mux2_1
XFILLER_192_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_255_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5789_ fd._0726_ fd._0894_ VGND VGND VPWR VPWR fd._0895_ sky130_fd_sc_hd__and2_1
XFILLER_130_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7528_ fd._2687_ VGND VGND VPWR VPWR fd._2808_ sky130_fd_sc_hd__clkinvlp_2
XTAP_5409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7459_ fd._2538_ fd._2731_ VGND VGND VPWR VPWR fd._2732_ sky130_fd_sc_hd__nand2_1
XTAP_4708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_1664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_268_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_279_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_273_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1559 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_231_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6830_ fd._2038_ fd._2039_ VGND VGND VPWR VPWR fd._2040_ sky130_fd_sc_hd__xnor2_1
XFILLER_19_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_208_ fd.c\[0\] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6761_ fd._1962_ fd._1963_ VGND VGND VPWR VPWR fd._1964_ sky130_fd_sc_hd__or2_1
XFILLER_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5712_ fd._0807_ fd._0809_ VGND VGND VPWR VPWR fd._0810_ sky130_fd_sc_hd__nand2_1
XFILLER_144_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6692_ fd._1645_ fd._1887_ VGND VGND VPWR VPWR fd._1888_ sky130_fd_sc_hd__nor2_1
XTAP_9270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5643_ fd._0568_ fd._0651_ VGND VGND VPWR VPWR fd._0734_ sky130_fd_sc_hd__or2_1
XFILLER_143_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._5574_ fd._0540_ fd._0657_ VGND VGND VPWR VPWR fd._0658_ sky130_fd_sc_hd__xnor2_1
XFILLER_174_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7313_ fd._2566_ fd._2570_ VGND VGND VPWR VPWR fd._2571_ sky130_fd_sc_hd__and2_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4525_ fd._3035_ fd._3598_ fd._3605_ VGND VGND VPWR VPWR fd._3619_ sky130_fd_sc_hd__o21ai_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7244_ fd._2492_ fd._2494_ VGND VGND VPWR VPWR fd._2495_ sky130_fd_sc_hd__nor2_1
XFILLER_22_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4456_ fd._2199_ fd._3387_ VGND VGND VPWR VPWR fd._3550_ sky130_fd_sc_hd__nor2_1
XFILLER_113_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_285_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_254_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_281_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7175_ fd._2325_ fd._2418_ VGND VGND VPWR VPWR fd._2420_ sky130_fd_sc_hd__xor2_1
XFILLER_93_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4387_ fd.b\[12\] fd._3416_ VGND VGND VPWR VPWR fd._3422_ sky130_fd_sc_hd__or2_1
XFILLER_226_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6126_ fd._1218_ fd._1225_ fd._1265_ fd._1226_ fd._1177_ VGND VGND VPWR VPWR fd._1266_
+ sky130_fd_sc_hd__o2111a_1
XFILLER_53_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_263_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._6057_ fd._1019_ VGND VGND VPWR VPWR fd._1190_ sky130_fd_sc_hd__clkinv_2
XFILLER_126_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5008_ fd._0025_ fd._0035_ fd._0033_ VGND VGND VPWR VPWR fd._0036_ sky130_fd_sc_hd__a21boi_1
XFILLER_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._6959_ fd._2169_ fd._2181_ VGND VGND VPWR VPWR fd._2182_ sky130_fd_sc_hd__or2b_1
XFILLER_162_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_260_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_268_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._4310_ fd.a\[15\] VGND VGND VPWR VPWR fd._2595_ sky130_fd_sc_hd__inv_2
XTAP_6496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5290_ fd._0345_ fd._0143_ VGND VGND VPWR VPWR fd._0346_ sky130_fd_sc_hd__xnor2_1
XFILLER_208_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_263_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4241_ fd._0219_ fd._1825_ VGND VGND VPWR VPWR fd._1836_ sky130_fd_sc_hd__xnor2_1
XFILLER_236_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4172_ fd._0835_ fd._0956_ fd._1066_ VGND VGND VPWR VPWR fd._1077_ sky130_fd_sc_hd__a21o_1
XFILLER_91_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_284_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7931_ fd._3223_ fd._3250_ VGND VGND VPWR VPWR fd._3251_ sky130_fd_sc_hd__xnor2_1
XFILLER_206_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7862_ fd._3163_ fd._3173_ fd._3174_ VGND VGND VPWR VPWR fd._3175_ sky130_fd_sc_hd__a21oi_1
XFILLER_15_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6813_ fd._1830_ fd._2019_ fd._2020_ VGND VGND VPWR VPWR fd._2021_ sky130_fd_sc_hd__mux2_1
XFILLER_121_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7793_ fd._1330_ fd._3098_ VGND VGND VPWR VPWR fd._3099_ sky130_fd_sc_hd__or2_1
XFILLER_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6744_ fd._1944_ fd._1936_ VGND VGND VPWR VPWR fd._1945_ sky130_fd_sc_hd__xnor2_1
XFILLER_89_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6675_ fd._1666_ fd._1868_ VGND VGND VPWR VPWR fd._1870_ sky130_fd_sc_hd__and2_1
XFILLER_144_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5626_ fd._3833_ VGND VGND VPWR VPWR fd._0716_ sky130_fd_sc_hd__buf_6
XFILLER_158_1592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_252_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_258_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5557_ fd._0262_ fd._0629_ fd._0636_ fd._0638_ fd._0639_ VGND VGND VPWR VPWR fd._0640_
+ sky130_fd_sc_hd__o221ai_2
XFILLER_119_1598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_273_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4508_ fd._3068_ fd._3601_ VGND VGND VPWR VPWR fd._3602_ sky130_fd_sc_hd__nand2_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_269_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5488_ fd._0555_ fd._0561_ fd._0563_ VGND VGND VPWR VPWR fd._0564_ sky130_fd_sc_hd__a21o_1
XFILLER_230_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_273_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_269_1554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7227_ fd._1816_ fd._2475_ VGND VGND VPWR VPWR fd._2477_ sky130_fd_sc_hd__nor2_1
XFILLER_38_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4439_ fd._3526_ fd._3532_ VGND VGND VPWR VPWR fd._3533_ sky130_fd_sc_hd__nand2_1
XFILLER_113_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7158_ fd._2206_ fd._2400_ VGND VGND VPWR VPWR fd._2401_ sky130_fd_sc_hd__xnor2_1
XFILLER_121_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6109_ fd._0716_ fd._1245_ VGND VGND VPWR VPWR fd._1247_ sky130_fd_sc_hd__nand2_1
XFILLER_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7089_ fd._1645_ fd._2324_ VGND VGND VPWR VPWR fd._2325_ sky130_fd_sc_hd__xnor2_1
XFILLER_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_263_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_277_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_249_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_242_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4790_ fd._3883_ fd._3860_ VGND VGND VPWR VPWR fd._3884_ sky130_fd_sc_hd__nor2_1
XFILLER_126_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6460_ fd._1434_ fd._1500_ fd._1502_ VGND VGND VPWR VPWR fd._1633_ sky130_fd_sc_hd__a21oi_1
XFILLER_206_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5411_ fd._3773_ VGND VGND VPWR VPWR fd._0479_ sky130_fd_sc_hd__buf_6
XFILLER_171_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6391_ fd._1555_ fd._1556_ VGND VGND VPWR VPWR fd._1557_ sky130_fd_sc_hd__or2_1
XTAP_6260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_255_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8130_ fd._3442_ fd._3443_ VGND VGND VPWR VPWR fd._3445_ sky130_fd_sc_hd__and2_1
XTAP_6282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_268_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5342_ fd._0200_ fd._0206_ fd._0209_ VGND VGND VPWR VPWR fd._0403_ sky130_fd_sc_hd__a21o_1
XTAP_6293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._8061_ fd._3364_ fd._3264_ fd._3386_ fd._3391_ fd._3393_ VGND VGND VPWR VPWR fd._3394_
+ sky130_fd_sc_hd__a311o_1
XFILLER_97_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5273_ fd._3675_ fd._0323_ VGND VGND VPWR VPWR fd._0327_ sky130_fd_sc_hd__or2_1
XFILLER_188_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_264_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7012_ fd._2235_ fd._2110_ VGND VGND VPWR VPWR fd._2240_ sky130_fd_sc_hd__nand2_1
XFILLER_75_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4224_ fd._0307_ fd._0406_ VGND VGND VPWR VPWR fd._1649_ sky130_fd_sc_hd__and2_1
XFILLER_224_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4155_ fd._0868_ fd.a\[10\] fd._0879_ fd._0604_ fd._0549_ VGND VGND VPWR VPWR
+ fd._0890_ sky130_fd_sc_hd__o221a_1
XFILLER_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_260_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4086_ fd.b\[19\] VGND VGND VPWR VPWR fd._0131_ sky130_fd_sc_hd__inv_6
XFILLER_176_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7914_ fd._3217_ fd._3052_ fd._3049_ VGND VGND VPWR VPWR fd._3232_ sky130_fd_sc_hd__o21a_1
XFILLER_31_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7845_ fd._3154_ fd._3155_ VGND VGND VPWR VPWR fd._3157_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._7776_ fd._2465_ fd._3078_ VGND VGND VPWR VPWR fd._3081_ sky130_fd_sc_hd__nor2_1
Xfd._4988_ fd._3580_ fd._0013_ VGND VGND VPWR VPWR fd._0014_ sky130_fd_sc_hd__nand2_1
XFILLER_118_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6727_ fd._1178_ fd._1743_ fd._1926_ VGND VGND VPWR VPWR fd._1927_ sky130_fd_sc_hd__a21o_1
XFILLER_160_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6658_ fd._1849_ fd._1850_ fd._1720_ VGND VGND VPWR VPWR fd._1851_ sky130_fd_sc_hd__mux2_1
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_263_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_258_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5609_ fd._0089_ fd._0694_ VGND VGND VPWR VPWR fd._0697_ sky130_fd_sc_hd__nor2_1
XFILLER_154_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6589_ fd._1559_ fd._1749_ VGND VGND VPWR VPWR fd._1775_ sky130_fd_sc_hd__or2_1
XFILLER_100_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_258_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8259_ net71 net11 VGND VGND VPWR VPWR fd.b\[19\] sky130_fd_sc_hd__dfxtp_2
XFILLER_227_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_254_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_1664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_1686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_250_1528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_283_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_261_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_261_1668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5960_ fd._0916_ fd._1082_ VGND VGND VPWR VPWR fd._1083_ sky130_fd_sc_hd__nor2_1
XFILLER_186_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4911_ fd._3869_ fd._4000_ fd._4004_ VGND VGND VPWR VPWR fd._4005_ sky130_fd_sc_hd__and3_1
XFILLER_224_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5891_ fd._0312_ fd._1006_ VGND VGND VPWR VPWR fd._1007_ sky130_fd_sc_hd__nor2_1
XFILLER_158_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7630_ fd._2912_ fd._2918_ fd._2919_ VGND VGND VPWR VPWR fd._2920_ sky130_fd_sc_hd__a21o_1
XFILLER_12_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4842_ fd._3795_ fd._3935_ VGND VGND VPWR VPWR fd._3936_ sky130_fd_sc_hd__nand2_1
Xuser_project_wrapper_100 VGND VGND VPWR VPWR user_project_wrapper_100/HI io_oeb[22]
+ sky130_fd_sc_hd__conb_1
XFILLER_220_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_project_wrapper_111 VGND VGND VPWR VPWR user_project_wrapper_111/HI io_oeb[33]
+ sky130_fd_sc_hd__conb_1
XFILLER_255_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_217_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_122 VGND VGND VPWR VPWR user_project_wrapper_122/HI la_data_out[0]
+ sky130_fd_sc_hd__conb_1
XFILLER_142_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7561_ fd._1242_ fd._2843_ VGND VGND VPWR VPWR fd._2844_ sky130_fd_sc_hd__nor2_1
Xuser_project_wrapper_133 VGND VGND VPWR VPWR user_project_wrapper_133/HI la_data_out[11]
+ sky130_fd_sc_hd__conb_1
Xfd._4773_ fd._3866_ fd._3686_ fd._3786_ VGND VGND VPWR VPWR fd._3867_ sky130_fd_sc_hd__mux2_1
XFILLER_182_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_144 VGND VGND VPWR VPWR user_project_wrapper_144/HI la_data_out[22]
+ sky130_fd_sc_hd__conb_1
XFILLER_5_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_255_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_project_wrapper_155 VGND VGND VPWR VPWR user_project_wrapper_155/HI la_data_out[33]
+ sky130_fd_sc_hd__conb_1
Xfd._6512_ fd._0965_ fd._1684_ fd._1689_ VGND VGND VPWR VPWR fd._1690_ sky130_fd_sc_hd__mux2_1
XFILLER_141_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_project_wrapper_166 VGND VGND VPWR VPWR user_project_wrapper_166/HI la_data_out[44]
+ sky130_fd_sc_hd__conb_1
XFILLER_99_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_177 VGND VGND VPWR VPWR user_project_wrapper_177/HI la_data_out[55]
+ sky130_fd_sc_hd__conb_1
Xfd._7492_ fd._2758_ fd._2764_ fd._2766_ fd._2767_ VGND VGND VPWR VPWR fd._2768_ sky130_fd_sc_hd__o31ai_2
XFILLER_138_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_project_wrapper_188 VGND VGND VPWR VPWR user_project_wrapper_188/HI la_data_out[66]
+ sky130_fd_sc_hd__conb_1
XFILLER_190_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_project_wrapper_199 VGND VGND VPWR VPWR user_project_wrapper_199/HI la_data_out[77]
+ sky130_fd_sc_hd__conb_1
XFILLER_218_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6443_ fd._1513_ fd._1524_ VGND VGND VPWR VPWR fd._1614_ sky130_fd_sc_hd__xor2_1
XFILLER_116_1524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_1415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_284_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_256_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_255_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6374_ fd._1405_ fd._1537_ VGND VGND VPWR VPWR fd._1538_ sky130_fd_sc_hd__xnor2_1
XFILLER_231_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8113_ fd._1231_ fd._3427_ VGND VGND VPWR VPWR fd._3428_ sky130_fd_sc_hd__nor2_1
XFILLER_256_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5325_ fd._0382_ fd._0383_ VGND VGND VPWR VPWR fd._0385_ sky130_fd_sc_hd__nor2_1
XFILLER_209_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8044_ fd._2465_ fd._3363_ fd._3374_ fd._2427_ VGND VGND VPWR VPWR fd._3375_ sky130_fd_sc_hd__o22a_1
Xfd._5256_ fd._3669_ fd._0308_ VGND VGND VPWR VPWR fd._0309_ sky130_fd_sc_hd__or2_1
XFILLER_3_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4207_ fd._0549_ VGND VGND VPWR VPWR fd._1462_ sky130_fd_sc_hd__inv_2
XFILLER_97_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5187_ fd._3947_ fd._0231_ VGND VGND VPWR VPWR fd._0233_ sky130_fd_sc_hd__nor2_2
XFILLER_211_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4138_ fd.a\[14\] fd.b\[14\] VGND VGND VPWR VPWR fd._0703_ sky130_fd_sc_hd__or2b_1
XFILLER_229_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_8409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7828_ fd._2929_ fd._3137_ VGND VGND VPWR VPWR fd._3138_ sky130_fd_sc_hd__xnor2_1
XFILLER_106_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7759_ fd._3021_ fd._3039_ fd._3051_ fd._3061_ VGND VGND VPWR VPWR fd._3062_ sky130_fd_sc_hd__o31a_1
XFILLER_106_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_259_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_275_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_274_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_261_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_265_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_265_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_230_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_8932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_269_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_266_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5110_ fd._0136_ fd._0140_ fd._0143_ fd._0144_ fd._0147_ VGND VGND VPWR VPWR fd._0148_
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_283_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6090_ fd._1219_ fd._1224_ VGND VGND VPWR VPWR fd._1226_ sky130_fd_sc_hd__nand2_1
XFILLER_19_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_283_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5041_ fd._0071_ VGND VGND VPWR VPWR fd._0072_ sky130_fd_sc_hd__clkinv_2
XTAP_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._6992_ fd._2002_ fd._2217_ fd._2116_ VGND VGND VPWR VPWR fd._2218_ sky130_fd_sc_hd__mux2_1
XFILLER_14_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._5943_ fd._0970_ fd._0973_ VGND VGND VPWR VPWR fd._1064_ sky130_fd_sc_hd__nor2_1
XFILLER_174_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5874_ fd._0839_ fd._0985_ fd._0986_ fd._0987_ VGND VGND VPWR VPWR fd._0988_ sky130_fd_sc_hd__o31a_1
XFILLER_31_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4825_ fd._3832_ fd._3918_ VGND VGND VPWR VPWR fd._3919_ sky130_fd_sc_hd__nand2_1
Xfd._7613_ fd._2773_ fd._2778_ fd._2781_ VGND VGND VPWR VPWR fd._2901_ sky130_fd_sc_hd__o21a_1
XFILLER_127_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_255_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4756_ fd._3849_ fd._3704_ fd._3787_ VGND VGND VPWR VPWR fd._3850_ sky130_fd_sc_hd__mux2_1
Xfd._7544_ fd._2645_ fd._2824_ VGND VGND VPWR VPWR fd._2825_ sky130_fd_sc_hd__and2_1
XFILLER_114_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_255_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7475_ fd._2142_ fd._2748_ VGND VGND VPWR VPWR fd._2750_ sky130_fd_sc_hd__or2_1
XFILLER_114_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4687_ fd._3767_ fd._3780_ VGND VGND VPWR VPWR fd._3781_ sky130_fd_sc_hd__and2b_1
XFILLER_151_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6426_ fd._1575_ fd._1593_ fd._1595_ fd._1573_ VGND VGND VPWR VPWR fd._1596_ sky130_fd_sc_hd__a211o_1
XFILLER_60_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_1578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6357_ fd._1313_ fd._1519_ fd._1423_ VGND VGND VPWR VPWR fd._1520_ sky130_fd_sc_hd__mux2_1
XFILLER_256_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_272_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5308_ fd._0364_ VGND VGND VPWR VPWR fd._0366_ sky130_fd_sc_hd__inv_2
XFILLER_37_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6288_ fd._0965_ fd._1443_ VGND VGND VPWR VPWR fd._1444_ sky130_fd_sc_hd__nand2_1
XFILLER_271_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8027_ fd._3351_ fd._3353_ fd._3341_ VGND VGND VPWR VPWR fd._3357_ sky130_fd_sc_hd__a21oi_1
XFILLER_37_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5239_ fd._0156_ fd._0289_ VGND VGND VPWR VPWR fd._0290_ sky130_fd_sc_hd__xnor2_1
XFILLER_164_1606 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_280_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_269_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_225_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_262_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_251_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_285_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_273_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_263_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_224_ fd.c\[16\] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_1
XFILLER_156_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_8751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4610_ fd._3507_ fd._3703_ fd._3624_ VGND VGND VPWR VPWR fd._3704_ sky130_fd_sc_hd__mux2_1
XFILLER_139_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._5590_ fd._0526_ fd._0675_ VGND VGND VPWR VPWR fd._0676_ sky130_fd_sc_hd__nand2_1
XFILLER_98_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4541_ fd._3629_ fd._3634_ VGND VGND VPWR VPWR fd._3635_ sky130_fd_sc_hd__nand2_1
XFILLER_151_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1690 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7260_ fd._2392_ fd._2498_ fd._2504_ VGND VGND VPWR VPWR fd._2513_ sky130_fd_sc_hd__and3_1
Xfd._4472_ fd._2562_ fd._2551_ VGND VGND VPWR VPWR fd._3566_ sky130_fd_sc_hd__and2b_1
XFILLER_239_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6211_ fd._0662_ fd._1358_ VGND VGND VPWR VPWR fd._1359_ sky130_fd_sc_hd__nor2_1
XFILLER_66_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7191_ fd._2274_ fd._2323_ VGND VGND VPWR VPWR fd._2437_ sky130_fd_sc_hd__nor2_1
XFILLER_120_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6142_ fd._1278_ fd._1281_ fd._1282_ VGND VGND VPWR VPWR fd._1283_ sky130_fd_sc_hd__o21ai_1
XFILLER_4_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_280_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6073_ fd._0632_ fd._1027_ VGND VGND VPWR VPWR fd._1207_ sky130_fd_sc_hd__nand2_1
XFILLER_280_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5024_ fd._0037_ VGND VGND VPWR VPWR fd._0053_ sky130_fd_sc_hd__inv_2
XFILLER_179_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6975_ fd._2196_ fd._2198_ fd._2115_ VGND VGND VPWR VPWR fd._2200_ sky130_fd_sc_hd__mux2_1
XFILLER_144_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5926_ fd._0998_ VGND VGND VPWR VPWR fd._1046_ sky130_fd_sc_hd__buf_6
XFILLER_175_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5857_ fd._0892_ fd._0969_ fd._0098_ VGND VGND VPWR VPWR fd._0970_ sky130_fd_sc_hd__o21a_1
XFILLER_179_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_274_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_255_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4808_ fd._3900_ fd._3901_ VGND VGND VPWR VPWR fd._3902_ sky130_fd_sc_hd__xnor2_1
Xfd._5788_ fd._0656_ fd._0893_ VGND VGND VPWR VPWR fd._0894_ sky130_fd_sc_hd__xnor2_1
XFILLER_157_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_255_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4739_ fd.b\[12\] VGND VGND VPWR VPWR fd._3833_ sky130_fd_sc_hd__buf_6
XFILLER_170_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7527_ fd._2698_ fd._2803_ fd._2806_ VGND VGND VPWR VPWR fd._2807_ sky130_fd_sc_hd__a21o_1
XFILLER_25_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_271_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7458_ fd._2533_ fd._2537_ VGND VGND VPWR VPWR fd._2731_ sky130_fd_sc_hd__or2_1
XTAP_4709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_272_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6409_ fd._0632_ fd._1399_ VGND VGND VPWR VPWR fd._1577_ sky130_fd_sc_hd__nor2_1
XFILLER_217_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7389_ fd._2465_ fd._2640_ VGND VGND VPWR VPWR fd._2655_ sky130_fd_sc_hd__nand2_1
XFILLER_268_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_257_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_281_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_262_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_1335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_267_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_1601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_262_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6760_ fd._1767_ fd._1960_ fd._1961_ VGND VGND VPWR VPWR fd._1963_ sky130_fd_sc_hd__a21oi_1
XFILLER_89_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5711_ fd._0622_ fd._0808_ fd._0801_ VGND VGND VPWR VPWR fd._0809_ sky130_fd_sc_hd__mux2_1
XFILLER_183_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6691_ fd._1863_ VGND VGND VPWR VPWR fd._1887_ sky130_fd_sc_hd__inv_2
XFILLER_128_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5642_ fd._0726_ fd._0569_ fd._0572_ VGND VGND VPWR VPWR fd._0733_ sky130_fd_sc_hd__o21ba_1
XTAP_9293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5573_ fd._0548_ fd._0547_ VGND VGND VPWR VPWR fd._0657_ sky130_fd_sc_hd__nor2_1
XFILLER_154_1638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4524_ fd._3613_ fd._3617_ VGND VGND VPWR VPWR fd._3618_ sky130_fd_sc_hd__nor2_1
XTAP_7891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7312_ fd._2567_ fd._2569_ fd._2505_ VGND VGND VPWR VPWR fd._2570_ sky130_fd_sc_hd__mux2_1
XFILLER_112_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._7243_ fd._1507_ fd._2493_ VGND VGND VPWR VPWR fd._2494_ sky130_fd_sc_hd__nor2_1
Xfd._4455_ fd._0428_ fd._3502_ fd._3545_ fd._3546_ fd._3548_ VGND VGND VPWR VPWR fd._3549_
+ sky130_fd_sc_hd__a2111o_1
XFILLER_254_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7174_ fd._2412_ fd._2416_ fd._2417_ VGND VGND VPWR VPWR fd._2418_ sky130_fd_sc_hd__a21oi_1
XFILLER_285_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4386_ fd._1561_ fd._3410_ fd._3211_ VGND VGND VPWR VPWR fd._3416_ sky130_fd_sc_hd__mux2_1
XFILLER_4_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6125_ fd._1262_ fd._1261_ VGND VGND VPWR VPWR fd._1265_ sky130_fd_sc_hd__and2b_1
XFILLER_0_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_1411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6056_ fd._0807_ fd._1188_ VGND VGND VPWR VPWR fd._1189_ sky130_fd_sc_hd__nand2_1
XFILLER_62_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5007_ fd._0033_ fd._0034_ VGND VGND VPWR VPWR fd._0035_ sky130_fd_sc_hd__and2_1
XFILLER_161_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_1628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6958_ fd._1585_ fd._1980_ VGND VGND VPWR VPWR fd._2181_ sky130_fd_sc_hd__nand2_1
XFILLER_175_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5909_ fd._0437_ fd._0858_ fd._0874_ fd._0984_ VGND VGND VPWR VPWR fd._1027_ sky130_fd_sc_hd__and4_1
XFILLER_107_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_266_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._6889_ fd._1304_ fd._2052_ VGND VGND VPWR VPWR fd._2105_ sky130_fd_sc_hd__nor2_1
XFILLER_190_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_249_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_244_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_285_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_281_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_257_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4240_ fd._1209_ fd._1792_ fd._1803_ fd._1814_ VGND VGND VPWR VPWR fd._1825_ sky130_fd_sc_hd__a31oi_2
XTAP_5796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_275_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4171_ fd._1000_ fd._1011_ fd._1022_ fd._1055_ VGND VGND VPWR VPWR fd._1066_ sky130_fd_sc_hd__or4b_1
XFILLER_78_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7930_ fd._3229_ fd._3227_ VGND VGND VPWR VPWR fd._3250_ sky130_fd_sc_hd__and2b_1
XFILLER_43_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7861_ fd._2142_ fd._3158_ VGND VGND VPWR VPWR fd._3174_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6812_ fd._1917_ VGND VGND VPWR VPWR fd._2020_ sky130_fd_sc_hd__buf_6
XFILLER_30_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7792_ fd._2996_ fd._3097_ fd._3076_ VGND VGND VPWR VPWR fd._3098_ sky130_fd_sc_hd__mux2_1
XFILLER_160_1697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6743_ fd._1774_ fd._1934_ VGND VGND VPWR VPWR fd._1944_ sky130_fd_sc_hd__and2_1
XFILLER_172_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6674_ fd._1648_ fd._1867_ fd._1720_ VGND VGND VPWR VPWR fd._1868_ sky130_fd_sc_hd__mux2_1
XFILLER_256_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5625_ fd._0712_ fd._0713_ VGND VGND VPWR VPWR fd._0715_ sky130_fd_sc_hd__or2_1
XFILLER_113_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5556_ fd._0125_ fd._0635_ fd._0631_ fd._0632_ VGND VGND VPWR VPWR fd._0639_ sky130_fd_sc_hd__a211o_1
XFILLER_113_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4507_ fd._3057_ fd._2969_ fd._3024_ VGND VGND VPWR VPWR fd._3601_ sky130_fd_sc_hd__nand3_1
XFILLER_239_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5487_ fd._0758_ fd._0562_ VGND VGND VPWR VPWR fd._0563_ sky130_fd_sc_hd__nor2_1
XFILLER_113_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4438_ fd.b\[0\] fd._3525_ VGND VGND VPWR VPWR fd._3532_ sky130_fd_sc_hd__nand2_1
Xfd._7226_ fd._1816_ fd._2475_ VGND VGND VPWR VPWR fd._2476_ sky130_fd_sc_hd__nand2_1
XFILLER_226_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4369_ fd._1440_ fd._2408_ VGND VGND VPWR VPWR fd._3244_ sky130_fd_sc_hd__nor2_1
XFILLER_226_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7157_ fd._1102_ fd._2211_ VGND VGND VPWR VPWR fd._2400_ sky130_fd_sc_hd__xnor2_1
XFILLER_148_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6108_ fd._0716_ fd._1245_ VGND VGND VPWR VPWR fd._1246_ sky130_fd_sc_hd__or2_1
Xfd._7088_ fd._2117_ fd._2230_ fd._2323_ VGND VGND VPWR VPWR fd._2324_ sky130_fd_sc_hd__mux2_1
XFILLER_223_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6039_ fd._0990_ fd._1039_ fd._1169_ VGND VGND VPWR VPWR fd._1170_ sky130_fd_sc_hd__mux2_1
XFILLER_22_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_260_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_268_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_267_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5410_ fd._0477_ fd._0460_ VGND VGND VPWR VPWR fd._0478_ sky130_fd_sc_hd__and2_2
XFILLER_150_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6390_ fd._1178_ fd._1554_ VGND VGND VPWR VPWR fd._1556_ sky130_fd_sc_hd__nor2_1
XFILLER_171_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5341_ fd._0401_ fd._0393_ VGND VGND VPWR VPWR fd._0402_ sky130_fd_sc_hd__and2_1
XFILLER_132_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_1643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._8060_ fd._3392_ fd._3262_ VGND VGND VPWR VPWR fd._3393_ sky130_fd_sc_hd__nor2_1
XFILLER_236_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5272_ fd._0312_ fd._0316_ VGND VGND VPWR VPWR fd._0326_ sky130_fd_sc_hd__nand2_1
XTAP_5593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4223_ fd.a\[5\] VGND VGND VPWR VPWR fd._1638_ sky130_fd_sc_hd__clkinv_2
Xfd._7011_ fd._2231_ fd._2237_ fd._2238_ VGND VGND VPWR VPWR fd._2239_ sky130_fd_sc_hd__mux2_1
XTAP_4881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._4154_ fd._0527_ VGND VGND VPWR VPWR fd._0879_ sky130_fd_sc_hd__inv_2
XFILLER_51_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4085_ fd._0065_ fd._0087_ fd._0109_ VGND VGND VPWR VPWR fd._0120_ sky130_fd_sc_hd__or3_1
XFILLER_264_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7913_ fd._3033_ VGND VGND VPWR VPWR fd._3231_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_203_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7844_ fd._2952_ fd._2961_ VGND VGND VPWR VPWR fd._3155_ sky130_fd_sc_hd__and2b_1
XFILLER_191_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7775_ fd._2465_ fd._3078_ VGND VGND VPWR VPWR fd._3080_ sky130_fd_sc_hd__nand2_1
Xfd._4987_ fd._3812_ fd._0012_ fd._3961_ VGND VGND VPWR VPWR fd._0013_ sky130_fd_sc_hd__mux2_1
XFILLER_69_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6726_ fd._1746_ fd._1750_ fd._1776_ VGND VGND VPWR VPWR fd._1926_ sky130_fd_sc_hd__nor3_1
XFILLER_144_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_275_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6657_ fd._1684_ fd._1689_ VGND VGND VPWR VPWR fd._1850_ sky130_fd_sc_hd__xnor2_1
XFILLER_160_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5608_ fd._0695_ VGND VGND VPWR VPWR fd._0696_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_258_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6588_ fd._1751_ fd._1755_ VGND VGND VPWR VPWR fd._1774_ sky130_fd_sc_hd__or2_1
XFILLER_113_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5539_ fd._0436_ fd._0619_ VGND VGND VPWR VPWR fd._0620_ sky130_fd_sc_hd__nand2_1
XFILLER_112_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_1590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8258_ net70 net10 VGND VGND VPWR VPWR fd.b\[18\] sky130_fd_sc_hd__dfxtp_2
XFILLER_269_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7209_ fd._2285_ fd._2456_ fd._2423_ VGND VGND VPWR VPWR fd._2457_ sky130_fd_sc_hd__mux2_1
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8189_ net72 fd.mc\[13\] VGND VGND VPWR VPWR fd.c\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_227_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_1601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_274_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4910_ fd._3954_ fd._3958_ fd._4003_ VGND VGND VPWR VPWR fd._4004_ sky130_fd_sc_hd__a21o_1
XFILLER_70_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5890_ fd._1005_ VGND VGND VPWR VPWR fd._1006_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_186_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4841_ fd._3803_ fd._3932_ fd._3934_ VGND VGND VPWR VPWR fd._3935_ sky130_fd_sc_hd__a21o_1
XFILLER_173_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_101 VGND VGND VPWR VPWR user_project_wrapper_101/HI io_oeb[23]
+ sky130_fd_sc_hd__conb_1
XFILLER_182_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_project_wrapper_112 VGND VGND VPWR VPWR user_project_wrapper_112/HI io_oeb[34]
+ sky130_fd_sc_hd__conb_1
XFILLER_103_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_project_wrapper_123 VGND VGND VPWR VPWR user_project_wrapper_123/HI la_data_out[1]
+ sky130_fd_sc_hd__conb_1
XFILLER_217_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7560_ fd._2635_ fd._2842_ fd._2813_ VGND VGND VPWR VPWR fd._2843_ sky130_fd_sc_hd__mux2_1
XFILLER_138_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4772_ fd._3863_ fd._3865_ VGND VGND VPWR VPWR fd._3866_ sky130_fd_sc_hd__xor2_1
XFILLER_126_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_134 VGND VGND VPWR VPWR user_project_wrapper_134/HI la_data_out[12]
+ sky130_fd_sc_hd__conb_1
XFILLER_99_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_145 VGND VGND VPWR VPWR user_project_wrapper_145/HI la_data_out[23]
+ sky130_fd_sc_hd__conb_1
XFILLER_5_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_156 VGND VGND VPWR VPWR user_project_wrapper_156/HI la_data_out[34]
+ sky130_fd_sc_hd__conb_1
XFILLER_177_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6511_ fd._1685_ fd._1688_ VGND VGND VPWR VPWR fd._1689_ sky130_fd_sc_hd__xnor2_1
Xuser_project_wrapper_167 VGND VGND VPWR VPWR user_project_wrapper_167/HI la_data_out[45]
+ sky130_fd_sc_hd__conb_1
XFILLER_29_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_178 VGND VGND VPWR VPWR user_project_wrapper_178/HI la_data_out[56]
+ sky130_fd_sc_hd__conb_1
XFILLER_269_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7491_ fd._2752_ fd._2757_ fd._2751_ VGND VGND VPWR VPWR fd._2767_ sky130_fd_sc_hd__a21o_1
XFILLER_99_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_189 VGND VGND VPWR VPWR user_project_wrapper_189/HI la_data_out[67]
+ sky130_fd_sc_hd__conb_1
XFILLER_116_1503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_269_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6442_ fd._1521_ VGND VGND VPWR VPWR fd._1613_ sky130_fd_sc_hd__clkinv_2
XFILLER_151_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_268_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6373_ fd._1536_ fd._1411_ VGND VGND VPWR VPWR fd._1537_ sky130_fd_sc_hd__nor2_1
XTAP_6080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_256_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8112_ fd._3425_ fd._3426_ VGND VGND VPWR VPWR fd._3427_ sky130_fd_sc_hd__nor2_1
XFILLER_231_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_284_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5324_ fd._0378_ VGND VGND VPWR VPWR fd._0383_ sky130_fd_sc_hd__inv_2
XFILLER_83_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_255_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5255_ fd._0103_ fd._0306_ fd._0268_ VGND VGND VPWR VPWR fd._0308_ sky130_fd_sc_hd__mux2_1
XFILLER_224_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._8043_ fd._3092_ fd._3241_ fd._3372_ fd._3373_ VGND VGND VPWR VPWR fd._3374_ sky130_fd_sc_hd__o22a_1
XFILLER_36_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_270_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4206_ fd.b\[12\] VGND VGND VPWR VPWR fd._1451_ sky130_fd_sc_hd__clkinv_4
XFILLER_149_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5186_ fd._3947_ fd._0231_ VGND VGND VPWR VPWR fd._0232_ sky130_fd_sc_hd__and2_1
XFILLER_52_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4137_ fd.b\[14\] fd.a\[14\] VGND VGND VPWR VPWR fd._0692_ sky130_fd_sc_hd__and2b_1
XFILLER_166_1670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7827_ fd._2934_ fd._2964_ VGND VGND VPWR VPWR fd._3137_ sky130_fd_sc_hd__nand2_1
XFILLER_69_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7758_ fd._3060_ VGND VGND VPWR VPWR fd._3061_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_69_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6709_ fd._0131_ fd._1906_ VGND VGND VPWR VPWR fd._1907_ sky130_fd_sc_hd__nor2_1
XFILLER_160_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_274_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7689_ fd._1872_ fd._2898_ VGND VGND VPWR VPWR fd._2985_ sky130_fd_sc_hd__nand2_1
XFILLER_121_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_243_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_243_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_284_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_283_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5040_ fd._4070_ fd._0006_ VGND VGND VPWR VPWR fd._0071_ sky130_fd_sc_hd__xor2_1
XFILLER_206_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_265_1591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._6991_ fd._2215_ fd._2216_ VGND VGND VPWR VPWR fd._2217_ sky130_fd_sc_hd__nor2_1
XFILLER_158_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5942_ fd._0877_ VGND VGND VPWR VPWR fd._1063_ sky130_fd_sc_hd__clkinv_2
XFILLER_13_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5873_ fd._0803_ fd._0985_ VGND VGND VPWR VPWR fd._0987_ sky130_fd_sc_hd__nand2_1
XFILLER_174_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7612_ fd._2717_ VGND VGND VPWR VPWR fd._2900_ sky130_fd_sc_hd__clkinv_2
XFILLER_122_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4824_ fd._3917_ fd._3831_ VGND VGND VPWR VPWR fd._3918_ sky130_fd_sc_hd__nand2_1
XFILLER_157_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7543_ fd._2427_ fd._2644_ VGND VGND VPWR VPWR fd._2824_ sky130_fd_sc_hd__nand2_1
XFILLER_138_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4755_ fd._3702_ fd._3848_ VGND VGND VPWR VPWR fd._3849_ sky130_fd_sc_hd__xnor2_1
XFILLER_103_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7474_ fd._2550_ fd._2747_ fd._2676_ VGND VGND VPWR VPWR fd._2748_ sky130_fd_sc_hd__mux2_1
Xfd._4686_ fd.b\[22\] fd._3766_ VGND VGND VPWR VPWR fd._3780_ sky130_fd_sc_hd__nand2_1
XFILLER_229_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6425_ fd._0807_ fd._1565_ VGND VGND VPWR VPWR fd._1595_ sky130_fd_sc_hd__nor2_1
XFILLER_68_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_256_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6356_ fd._1518_ VGND VGND VPWR VPWR fd._1519_ sky130_fd_sc_hd__clkinv_2
XFILLER_3_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5307_ fd._0758_ fd._0364_ VGND VGND VPWR VPWR fd._0365_ sky130_fd_sc_hd__nor2_1
XFILLER_209_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6287_ fd._1288_ fd._1442_ fd._1422_ VGND VGND VPWR VPWR fd._1443_ sky130_fd_sc_hd__mux2_1
XFILLER_37_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8026_ fd._3307_ fd._3308_ fd._3322_ fd._3333_ fd._3355_ VGND VGND VPWR VPWR fd._3356_
+ sky130_fd_sc_hd__a2111oi_2
XFILLER_77_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5238_ fd._0163_ fd._0162_ VGND VGND VPWR VPWR fd._0289_ sky130_fd_sc_hd__or2b_1
XFILLER_225_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1618 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_251_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5169_ fd._0016_ fd._0212_ VGND VGND VPWR VPWR fd._0213_ sky130_fd_sc_hd__xnor2_1
XFILLER_24_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_269_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_1517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_225_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_1686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_279_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_273_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_273_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_266_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_259_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_275_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_256_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_243_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_223_ fd.c\[15\] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_1
XFILLER_230_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_256_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4540_ fd._3565_ fd._3569_ VGND VGND VPWR VPWR fd._3634_ sky130_fd_sc_hd__or2_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4471_ fd._3332_ fd._3459_ fd._3564_ VGND VGND VPWR VPWR fd._3565_ sky130_fd_sc_hd__or3_1
XFILLER_214_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6210_ fd._1357_ VGND VGND VPWR VPWR fd._1358_ sky130_fd_sc_hd__inv_2
XFILLER_254_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._7190_ fd._2270_ fd._2435_ VGND VGND VPWR VPWR fd._2436_ sky130_fd_sc_hd__xnor2_1
XFILLER_66_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6141_ fd._0726_ fd._1240_ VGND VGND VPWR VPWR fd._1282_ sky130_fd_sc_hd__nand2_1
XFILLER_92_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6072_ fd._3695_ fd._1059_ fd._1074_ fd._1167_ VGND VGND VPWR VPWR fd._1206_ sky130_fd_sc_hd__or4_2
XFILLER_74_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5023_ fd._0037_ fd._0033_ fd._0051_ fd._3967_ VGND VGND VPWR VPWR fd._0052_ sky130_fd_sc_hd__a211o_1
XFILLER_228_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6974_ fd._1996_ fd._2197_ VGND VGND VPWR VPWR fd._2198_ sky130_fd_sc_hd__xor2_1
XFILLER_72_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5925_ fd._1043_ VGND VGND VPWR VPWR fd._1045_ sky130_fd_sc_hd__clkinv_2
XFILLER_119_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5856_ fd._0960_ fd._0964_ fd._0966_ fd._0968_ VGND VGND VPWR VPWR fd._0969_ sky130_fd_sc_hd__o211a_1
XFILLER_161_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_255_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_255_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4807_ fd._3714_ fd._3654_ VGND VGND VPWR VPWR fd._3901_ sky130_fd_sc_hd__nor2_1
XFILLER_161_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5787_ fd._0723_ fd._0722_ fd._0848_ VGND VGND VPWR VPWR fd._0893_ sky130_fd_sc_hd__nand3b_1
XFILLER_118_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7526_ fd._2805_ VGND VGND VPWR VPWR fd._2806_ sky130_fd_sc_hd__clkinv_4
XFILLER_255_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4738_ fd.b\[13\] fd._3831_ VGND VGND VPWR VPWR fd._3832_ sky130_fd_sc_hd__or2_1
XFILLER_130_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_257_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7457_ fd._2544_ fd._2552_ fd._2558_ fd._2559_ VGND VGND VPWR VPWR fd._2730_ sky130_fd_sc_hd__a31o_1
XFILLER_124_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4669_ fd._3760_ fd._3762_ fd._3626_ VGND VGND VPWR VPWR fd._3763_ sky130_fd_sc_hd__mux2_1
XFILLER_130_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6408_ fd._1393_ fd._1395_ VGND VGND VPWR VPWR fd._1576_ sky130_fd_sc_hd__or2_1
XFILLER_112_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_256_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7388_ fd._2427_ fd._2644_ fd._2646_ fd._2652_ fd._2653_ VGND VGND VPWR VPWR fd._2654_
+ sky130_fd_sc_hd__a221o_1
XFILLER_272_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6339_ fd._1438_ fd._1496_ fd._1498_ fd._1499_ VGND VGND VPWR VPWR fd._1500_ sky130_fd_sc_hd__a211o_1
XFILLER_17_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_272_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_281_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_262_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8009_ fd._3109_ fd._3336_ fd._3240_ VGND VGND VPWR VPWR fd._3337_ sky130_fd_sc_hd__mux2_1
XFILLER_266_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_262_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_240_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_8059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_1563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_251_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_249_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_284_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_280_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1550 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_28 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._5710_ fd._0623_ fd._0641_ VGND VGND VPWR VPWR fd._0808_ sky130_fd_sc_hd__xnor2_1
XFILLER_156_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6690_ fd._1879_ fd._1884_ fd._1885_ VGND VGND VPWR VPWR fd._1886_ sky130_fd_sc_hd__a21bo_1
XFILLER_32_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_9261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5641_ fd._0726_ fd._0564_ fd._0568_ VGND VGND VPWR VPWR fd._0732_ sky130_fd_sc_hd__and3_1
XFILLER_143_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5572_ fd._0654_ fd._0655_ fd._0651_ VGND VGND VPWR VPWR fd._0656_ sky130_fd_sc_hd__mux2_1
XFILLER_112_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7311_ fd._2396_ fd._2568_ VGND VGND VPWR VPWR fd._2569_ sky130_fd_sc_hd__xnor2_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4523_ fd._3614_ fd._3616_ fd._3222_ VGND VGND VPWR VPWR fd._3617_ sky130_fd_sc_hd__mux2_1
XFILLER_239_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_285_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_1674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7242_ fd._2491_ VGND VGND VPWR VPWR fd._2493_ sky130_fd_sc_hd__inv_2
Xfd._4454_ fd._3496_ fd._3547_ VGND VGND VPWR VPWR fd._3548_ sky130_fd_sc_hd__nand2_1
XFILLER_113_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7173_ fd._2093_ fd._2415_ VGND VGND VPWR VPWR fd._2417_ sky130_fd_sc_hd__nor2_1
XFILLER_113_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4385_ fd._2331_ fd._3404_ VGND VGND VPWR VPWR fd._3410_ sky130_fd_sc_hd__xnor2_1
XFILLER_253_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_254_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_285_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6124_ fd._1261_ fd._1174_ fd._1262_ VGND VGND VPWR VPWR fd._1263_ sky130_fd_sc_hd__a21oi_1
XFILLER_4_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_263_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6055_ fd._1013_ fd._1186_ fd._1169_ VGND VGND VPWR VPWR fd._1188_ sky130_fd_sc_hd__mux2_1
XFILLER_59_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5006_ fd._0026_ fd._0031_ VGND VGND VPWR VPWR fd._0034_ sky130_fd_sc_hd__nand2_1
XFILLER_210_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6957_ fd._1970_ fd._2020_ VGND VGND VPWR VPWR fd._2180_ sky130_fd_sc_hd__nand2_1
XFILLER_120_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5908_ fd._0858_ fd._0874_ fd._0984_ fd._1023_ VGND VGND VPWR VPWR fd._1026_ sky130_fd_sc_hd__a31o_1
XFILLER_175_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6888_ fd._2075_ fd._2102_ fd._2103_ fd._2073_ VGND VGND VPWR VPWR fd._2104_ sky130_fd_sc_hd__o211a_1
XFILLER_274_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._5839_ fd._0541_ fd._0946_ VGND VGND VPWR VPWR fd._0950_ sky130_fd_sc_hd__nand2_1
XFILLER_200_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_249_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7509_ fd._2570_ VGND VGND VPWR VPWR fd._2787_ sky130_fd_sc_hd__clkinv_2
XFILLER_130_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_268_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_257_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_272_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_260_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_281_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_281_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_268_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_268_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_267_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4170_ fd._0087_ fd._1044_ VGND VGND VPWR VPWR fd._1055_ sky130_fd_sc_hd__nor2_1
XFILLER_229_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_251_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7860_ fd._2751_ fd._3162_ fd._3169_ fd._3171_ fd._3172_ VGND VGND VPWR VPWR fd._3173_
+ sky130_fd_sc_hd__a221o_1
XFILLER_15_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6811_ fd._2018_ fd._1832_ VGND VGND VPWR VPWR fd._2019_ sky130_fd_sc_hd__xnor2_1
XFILLER_15_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7791_ fd._2997_ fd._2992_ VGND VGND VPWR VPWR fd._3097_ sky130_fd_sc_hd__xnor2_1
XFILLER_89_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_258_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6742_ fd._1941_ fd._1942_ VGND VGND VPWR VPWR fd._1943_ sky130_fd_sc_hd__nand2_1
XFILLER_157_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6673_ fd._1659_ fd._1662_ fd._1865_ fd._1866_ VGND VGND VPWR VPWR fd._1867_ sky130_fd_sc_hd__a31o_1
XFILLER_176_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_256_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5624_ fd._0541_ fd._0711_ VGND VGND VPWR VPWR fd._0713_ sky130_fd_sc_hd__nor2_1
XFILLER_193_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_8390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_271_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5555_ fd._0125_ VGND VGND VPWR VPWR fd._0638_ sky130_fd_sc_hd__buf_6
XFILLER_113_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4506_ fd._3592_ fd._3594_ fd._3599_ VGND VGND VPWR VPWR fd._3600_ sky130_fd_sc_hd__a21oi_2
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_252_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5486_ fd._0559_ VGND VGND VPWR VPWR fd._0562_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_22_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7225_ fd._2311_ fd._2473_ fd._2423_ VGND VGND VPWR VPWR fd._2475_ sky130_fd_sc_hd__mux2_1
XFILLER_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4437_ fd.b\[3\] fd._3530_ VGND VGND VPWR VPWR fd._3531_ sky130_fd_sc_hd__and2_1
XFILLER_22_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7156_ fd._2335_ fd._2347_ fd._2398_ fd._2333_ VGND VGND VPWR VPWR fd._2399_ sky130_fd_sc_hd__o31a_1
XFILLER_54_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_282_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4368_ fd._1374_ fd._2727_ fd._3222_ VGND VGND VPWR VPWR fd._3233_ sky130_fd_sc_hd__mux2_1
XFILLER_199_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6107_ fd._1108_ fd._1244_ fd._1223_ VGND VGND VPWR VPWR fd._1245_ sky130_fd_sc_hd__mux2_1
XFILLER_187_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7087_ fd._2322_ VGND VGND VPWR VPWR fd._2323_ sky130_fd_sc_hd__buf_6
XFILLER_53_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4299_ fd.b\[14\] fd._2452_ VGND VGND VPWR VPWR fd._2474_ sky130_fd_sc_hd__or2_1
XFILLER_263_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6038_ fd._1168_ VGND VGND VPWR VPWR fd._1169_ sky130_fd_sc_hd__buf_6
XFILLER_224_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_263_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7989_ fd._3135_ fd._3314_ fd._3132_ VGND VGND VPWR VPWR fd._3315_ sky130_fd_sc_hd__a21o_1
XFILLER_241_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1672 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_258_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1618 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5340_ fd._1352_ fd._0400_ VGND VGND VPWR VPWR fd._0401_ sky130_fd_sc_hd__or2_1
XTAP_6273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5271_ fd._0261_ fd._0257_ fd._0259_ fd._0264_ VGND VGND VPWR VPWR fd._0325_ sky130_fd_sc_hd__o31a_1
XTAP_5583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7010_ fd._2116_ VGND VGND VPWR VPWR fd._2238_ sky130_fd_sc_hd__clkbuf_4
XTAP_4871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4222_ fd._0857_ fd._1583_ fd._1605_ fd._1616_ VGND VGND VPWR VPWR fd._1627_ sky130_fd_sc_hd__o31a_1
XFILLER_188_1554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4153_ fd._0857_ VGND VGND VPWR VPWR fd._0868_ sky130_fd_sc_hd__clkinv_2
XFILLER_223_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4084_ fd._0098_ fd.a\[17\] VGND VGND VPWR VPWR fd._0109_ sky130_fd_sc_hd__nor2_1
XFILLER_189_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7912_ fd._3223_ fd._3227_ fd._3228_ fd._3229_ VGND VGND VPWR VPWR fd._3230_ sky130_fd_sc_hd__a211o_1
XFILLER_231_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7843_ fd._2957_ fd._2960_ VGND VGND VPWR VPWR fd._3154_ sky130_fd_sc_hd__or2_1
XFILLER_34_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7774_ fd._3070_ fd._3072_ fd._3077_ VGND VGND VPWR VPWR fd._3078_ sky130_fd_sc_hd__mux2_1
XFILLER_121_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._4986_ fd._0009_ fd._0011_ VGND VGND VPWR VPWR fd._0012_ sky130_fd_sc_hd__xnor2_1
XFILLER_247_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6725_ fd._1600_ fd._1923_ VGND VGND VPWR VPWR fd._1925_ sky130_fd_sc_hd__or2_1
XFILLER_105_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6656_ fd._1688_ VGND VGND VPWR VPWR fd._1849_ sky130_fd_sc_hd__clkinv_2
XFILLER_28_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_275_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._5607_ fd._0089_ fd._0694_ VGND VGND VPWR VPWR fd._0695_ sky130_fd_sc_hd__nand2_1
XFILLER_113_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6587_ fd._1015_ fd._1761_ fd._1767_ fd._1772_ VGND VGND VPWR VPWR fd._1773_ sky130_fd_sc_hd__o211a_1
XFILLER_112_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5538_ fd._0262_ fd._0435_ VGND VGND VPWR VPWR fd._0619_ sky130_fd_sc_hd__or2_1
XFILLER_171_1580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_258_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8257_ net70 net9 VGND VGND VPWR VPWR fd.b\[17\] sky130_fd_sc_hd__dfxtp_2
XFILLER_273_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5469_ fd._0303_ fd._0342_ VGND VGND VPWR VPWR fd._0543_ sky130_fd_sc_hd__nand2_1
XFILLER_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_269_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7208_ fd._1685_ fd._2455_ VGND VGND VPWR VPWR fd._2456_ sky130_fd_sc_hd__xnor2_1
XFILLER_132_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8188_ net74 fd.mc\[12\] VGND VGND VPWR VPWR fd.c\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_167_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_242_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_282_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7139_ fd._2376_ fd._2379_ fd._1976_ VGND VGND VPWR VPWR fd._2380_ sky130_fd_sc_hd__o21ai_1
XFILLER_148_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_282_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_1431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1032 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_1390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4840_ fd._3795_ fd._3933_ VGND VGND VPWR VPWR fd._3934_ sky130_fd_sc_hd__nand2_1
XFILLER_31_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_102 VGND VGND VPWR VPWR user_project_wrapper_102/HI io_oeb[24]
+ sky130_fd_sc_hd__conb_1
XFILLER_177_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_113 VGND VGND VPWR VPWR user_project_wrapper_113/HI io_oeb[35]
+ sky130_fd_sc_hd__conb_1
Xfd._4771_ fd._3687_ fd._3864_ VGND VGND VPWR VPWR fd._3865_ sky130_fd_sc_hd__nand2_1
Xuser_project_wrapper_124 VGND VGND VPWR VPWR user_project_wrapper_124/HI la_data_out[2]
+ sky130_fd_sc_hd__conb_1
XFILLER_192_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xuser_project_wrapper_135 VGND VGND VPWR VPWR user_project_wrapper_135/HI la_data_out[13]
+ sky130_fd_sc_hd__conb_1
XFILLER_259_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_146 VGND VGND VPWR VPWR user_project_wrapper_146/HI la_data_out[24]
+ sky130_fd_sc_hd__conb_1
XFILLER_86_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6510_ fd._1487_ fd._1687_ fd._1615_ VGND VGND VPWR VPWR fd._1688_ sky130_fd_sc_hd__mux2_1
XFILLER_126_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_157 VGND VGND VPWR VPWR user_project_wrapper_157/HI la_data_out[35]
+ sky130_fd_sc_hd__conb_1
XFILLER_5_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7490_ fd._1976_ fd._2759_ fd._2762_ fd._2377_ fd._2765_ VGND VGND VPWR VPWR fd._2766_
+ sky130_fd_sc_hd__o32a_1
Xuser_project_wrapper_168 VGND VGND VPWR VPWR user_project_wrapper_168/HI la_data_out[46]
+ sky130_fd_sc_hd__conb_1
XFILLER_253_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_179 VGND VGND VPWR VPWR user_project_wrapper_179/HI la_data_out[57]
+ sky130_fd_sc_hd__conb_1
XFILLER_269_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_268_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6441_ fd._1608_ fd._1611_ VGND VGND VPWR VPWR fd._1612_ sky130_fd_sc_hd__xnor2_1
XFILLER_214_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_284_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6372_ fd._0928_ fd._1409_ VGND VGND VPWR VPWR fd._1536_ sky130_fd_sc_hd__nor2_1
XTAP_6070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._8111_ fd.a\[23\] fd.b\[23\] VGND VGND VPWR VPWR fd._3426_ sky130_fd_sc_hd__and2b_1
XTAP_6092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5323_ fd._1308_ VGND VGND VPWR VPWR fd._0382_ sky130_fd_sc_hd__clkinv_4
XFILLER_255_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_1504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._8042_ fd._3370_ fd._3371_ fd._3241_ VGND VGND VPWR VPWR fd._3373_ sky130_fd_sc_hd__a21bo_1
XFILLER_76_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_252_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5254_ fd._0304_ fd._0305_ VGND VGND VPWR VPWR fd._0306_ sky130_fd_sc_hd__xor2_1
XFILLER_23_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_264_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4205_ fd.b\[13\] fd._1429_ VGND VGND VPWR VPWR fd._1440_ sky130_fd_sc_hd__nor2_1
XFILLER_188_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_263_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5185_ fd._3966_ fd._0229_ fd._0061_ VGND VGND VPWR VPWR fd._0231_ sky130_fd_sc_hd__mux2_1
XFILLER_224_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4136_ fd._0659_ fd._0670_ VGND VGND VPWR VPWR fd._0681_ sky130_fd_sc_hd__and2b_1
XFILLER_166_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_264_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7826_ fd._3135_ VGND VGND VPWR VPWR fd._3136_ sky130_fd_sc_hd__inv_2
XFILLER_157_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7757_ fd._3049_ fd._3038_ fd._3052_ fd._3059_ VGND VGND VPWR VPWR fd._3060_ sky130_fd_sc_hd__a31o_1
XFILLER_121_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4969_ fd._4063_ fd._4064_ VGND VGND VPWR VPWR fd._4065_ sky130_fd_sc_hd__xor2_1
XFILLER_160_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6708_ fd._1841_ VGND VGND VPWR VPWR fd._1906_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_145_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7688_ fd._1656_ fd._2983_ VGND VGND VPWR VPWR fd._2984_ sky130_fd_sc_hd__nand2_1
XFILLER_47_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6639_ fd._1819_ VGND VGND VPWR VPWR fd._1830_ sky130_fd_sc_hd__inv_2
XFILLER_8_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_255_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_1643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_8967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_1583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_266_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_261_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_1576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6990_ fd._1933_ fd._1997_ fd._2214_ VGND VGND VPWR VPWR fd._2216_ sky130_fd_sc_hd__a21oi_1
XFILLER_20_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5941_ fd._0479_ fd._1061_ VGND VGND VPWR VPWR fd._1062_ sky130_fd_sc_hd__nor2_1
XFILLER_201_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5872_ fd._0810_ fd._0838_ fd._0806_ VGND VGND VPWR VPWR fd._0986_ sky130_fd_sc_hd__a21oi_1
XFILLER_179_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7611_ fd._1872_ fd._2898_ VGND VGND VPWR VPWR fd._2899_ sky130_fd_sc_hd__or2_1
Xfd._4823_ fd.b\[13\] VGND VGND VPWR VPWR fd._3917_ sky130_fd_sc_hd__buf_6
XFILLER_196_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7542_ fd._2646_ fd._2652_ fd._2653_ VGND VGND VPWR VPWR fd._2823_ sky130_fd_sc_hd__a21oi_1
XFILLER_127_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4754_ fd._3709_ fd._3705_ VGND VGND VPWR VPWR fd._3848_ sky130_fd_sc_hd__or2b_1
XFILLER_192_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_269_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7473_ fd._2744_ fd._2746_ VGND VGND VPWR VPWR fd._2747_ sky130_fd_sc_hd__xnor2_1
Xfd._4685_ fd._3035_ fd._3755_ fd._3778_ VGND VGND VPWR VPWR fd._3779_ sky130_fd_sc_hd__o21a_1
XFILLER_155_1350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6424_ fd._1582_ fd._1589_ fd._1591_ fd._1592_ VGND VGND VPWR VPWR fd._1593_ sky130_fd_sc_hd__o31ai_2
XFILLER_269_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_256_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6355_ fd._1316_ fd._1516_ VGND VGND VPWR VPWR fd._1518_ sky130_fd_sc_hd__xnor2_1
XFILLER_151_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_249_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5306_ fd._0079_ fd._0363_ fd._0269_ VGND VGND VPWR VPWR fd._0364_ sky130_fd_sc_hd__mux2_1
XFILLER_83_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6286_ fd._1439_ fd._1441_ VGND VGND VPWR VPWR fd._1442_ sky130_fd_sc_hd__xnor2_1
XFILLER_114_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8025_ fd._3341_ fd._3342_ fd._3352_ fd._3353_ VGND VGND VPWR VPWR fd._3355_ sky130_fd_sc_hd__or4bb_1
Xfd._5237_ fd._0000_ fd._0287_ VGND VGND VPWR VPWR fd._0288_ sky130_fd_sc_hd__or2_1
XFILLER_36_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5168_ fd._0024_ fd._0023_ VGND VGND VPWR VPWR fd._0212_ sky130_fd_sc_hd__or2b_1
XFILLER_52_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4119_ fd.b\[7\] fd._0439_ fd.b\[6\] fd._0483_ VGND VGND VPWR VPWR fd._0494_ sky130_fd_sc_hd__a211o_1
XFILLER_240_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_264_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_1676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5099_ fd._0100_ fd._0105_ fd._0135_ fd._0097_ VGND VGND VPWR VPWR fd._0136_ sky130_fd_sc_hd__a31o_1
XFILLER_127_1496 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_8219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7809_ fd._3111_ fd._3116_ VGND VGND VPWR VPWR fd._3117_ sky130_fd_sc_hd__nor2_1
XFILLER_192_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_251_1658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_219_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_284_1412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_227_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_222_ fd.c\[14\] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_1
XFILLER_243_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4470_ fd._3555_ fd._3558_ fd._3563_ VGND VGND VPWR VPWR fd._3564_ sky130_fd_sc_hd__a21oi_1
XFILLER_6_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_1580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6140_ fd._1118_ fd._1277_ fd._1280_ VGND VGND VPWR VPWR fd._1281_ sky130_fd_sc_hd__a21oi_1
XFILLER_65_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_219_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6071_ fd._0318_ fd._1204_ VGND VGND VPWR VPWR fd._1205_ sky130_fd_sc_hd__or2_1
XFILLER_18_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5022_ fd._0046_ fd._0041_ VGND VGND VPWR VPWR fd._0051_ sky130_fd_sc_hd__or2_1
XFILLER_206_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_261_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._6973_ fd._1986_ fd._1991_ fd._1994_ VGND VGND VPWR VPWR fd._2197_ sky130_fd_sc_hd__a21oi_1
XFILLER_261_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5924_ fd._1042_ fd._0872_ VGND VGND VPWR VPWR fd._1043_ sky130_fd_sc_hd__xor2_1
XFILLER_105_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_1502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5855_ fd._1308_ fd._0963_ VGND VGND VPWR VPWR fd._0968_ sky130_fd_sc_hd__nand2_1
XFILLER_134_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4806_ fd._3663_ fd._3710_ VGND VGND VPWR VPWR fd._3900_ sky130_fd_sc_hd__nand2_1
XFILLER_255_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5786_ fd._0891_ VGND VGND VPWR VPWR fd._0892_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_143_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_255_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7525_ fd._1330_ fd._2691_ VGND VGND VPWR VPWR fd._2805_ sky130_fd_sc_hd__xnor2_1
Xfd._4737_ fd._3829_ fd._3788_ fd._3830_ VGND VGND VPWR VPWR fd._3831_ sky130_fd_sc_hd__o21a_1
XFILLER_153_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7456_ fd._2537_ VGND VGND VPWR VPWR fd._2729_ sky130_fd_sc_hd__clkinv_2
Xfd._4668_ fd._3613_ fd._3761_ VGND VGND VPWR VPWR fd._3762_ sky130_fd_sc_hd__xnor2_1
XFILLER_124_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_256_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6407_ fd._1573_ fd._1574_ VGND VGND VPWR VPWR fd._1575_ sky130_fd_sc_hd__nor2b_1
XFILLER_271_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7387_ fd._1286_ fd._2651_ VGND VGND VPWR VPWR fd._2653_ sky130_fd_sc_hd__and2_1
XFILLER_84_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4599_ fd._3690_ fd._3692_ fd._3624_ VGND VGND VPWR VPWR fd._3693_ sky130_fd_sc_hd__mux2_1
XFILLER_112_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_268_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_256_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6338_ fd._0098_ fd._1444_ fd._1493_ VGND VGND VPWR VPWR fd._1499_ sky130_fd_sc_hd__and3_1
XFILLER_68_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6269_ fd._1422_ VGND VGND VPWR VPWR fd._1423_ sky130_fd_sc_hd__buf_6
XFILLER_168_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8008_ fd._3335_ fd._3201_ VGND VGND VPWR VPWR fd._3336_ sky130_fd_sc_hd__xor2_1
XFILLER_77_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_266_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_1560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_279_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_273_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_273_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_251_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_1575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_250_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_249_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_262_1562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5640_ fd._0724_ fd._0726_ fd._0730_ VGND VGND VPWR VPWR fd._0731_ sky130_fd_sc_hd__mux2_1
XFILLER_193_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5571_ fd._0550_ fd._0554_ VGND VGND VPWR VPWR fd._0655_ sky130_fd_sc_hd__xnor2_1
XFILLER_140_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_285_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7310_ fd._2389_ fd._2393_ fd._2395_ VGND VGND VPWR VPWR fd._2568_ sky130_fd_sc_hd__o21a_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4522_ fd._3134_ fd._3615_ VGND VGND VPWR VPWR fd._3616_ sky130_fd_sc_hd__xnor2_1
XTAP_7871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_285_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7241_ fd._1242_ fd._2491_ VGND VGND VPWR VPWR fd._2492_ sky130_fd_sc_hd__nor2_1
XFILLER_269_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4453_ fd._2155_ fd._3495_ VGND VGND VPWR VPWR fd._3547_ sky130_fd_sc_hd__nand2_1
XFILLER_234_1697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_254_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7172_ fd._2093_ fd._2415_ VGND VGND VPWR VPWR fd._2416_ sky130_fd_sc_hd__nand2_1
XFILLER_43_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4384_ fd._3397_ fd._2342_ fd._0857_ fd._1605_ VGND VGND VPWR VPWR fd._3404_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_130_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6123_ fd._0916_ fd._1260_ VGND VGND VPWR VPWR fd._1262_ sky130_fd_sc_hd__and2_1
XFILLER_24_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_254_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_267_1484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6054_ fd._1014_ fd._1179_ VGND VGND VPWR VPWR fd._1186_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5005_ fd._0026_ fd._0031_ VGND VGND VPWR VPWR fd._0033_ sky130_fd_sc_hd__or2_1
XFILLER_206_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_1668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6956_ fd._2175_ fd._2176_ fd._2178_ VGND VGND VPWR VPWR fd._2179_ sky130_fd_sc_hd__and3_1
XFILLER_30_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5907_ fd._0985_ fd._1021_ fd._1024_ fd._0638_ VGND VGND VPWR VPWR fd._1025_ sky130_fd_sc_hd__a211o_1
XFILLER_190_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6887_ fd._1275_ fd._2065_ VGND VGND VPWR VPWR fd._2103_ sky130_fd_sc_hd__nand2_1
XFILLER_135_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5838_ fd._0903_ fd._0948_ VGND VGND VPWR VPWR fd._0949_ sky130_fd_sc_hd__nand2_1
XFILLER_157_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5769_ fd._0850_ fd._0872_ VGND VGND VPWR VPWR fd._0873_ sky130_fd_sc_hd__nor2_1
XFILLER_130_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7508_ fd._2773_ fd._2778_ fd._2779_ fd._2781_ fd._2785_ VGND VGND VPWR VPWR fd._2786_
+ sky130_fd_sc_hd__o2111a_1
XFILLER_118_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_257_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7439_ fd._1797_ fd._2709_ VGND VGND VPWR VPWR fd._2710_ sky130_fd_sc_hd__and2_1
XFILLER_28_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_257_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_268_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_275_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_284_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_262_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_231_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6810_ fd._1824_ fd._2017_ fd._1834_ VGND VGND VPWR VPWR fd._2018_ sky130_fd_sc_hd__a21o_1
XFILLER_200_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7790_ fd._1685_ fd._3095_ VGND VGND VPWR VPWR fd._3096_ sky130_fd_sc_hd__nand2_1
XFILLER_15_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6741_ fd._0504_ fd._1940_ VGND VGND VPWR VPWR fd._1942_ sky130_fd_sc_hd__nand2_1
XFILLER_172_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6672_ fd._0716_ fd._1659_ VGND VGND VPWR VPWR fd._1866_ sky130_fd_sc_hd__nor2_1
XTAP_9070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5623_ fd._0541_ fd._0711_ VGND VGND VPWR VPWR fd._0712_ sky130_fd_sc_hd__and2_1
XFILLER_119_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_259_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_252_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5554_ fd._0453_ fd._0631_ fd._0635_ VGND VGND VPWR VPWR fd._0636_ sky130_fd_sc_hd__a21boi_2
XFILLER_140_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4505_ fd._3035_ fd._3598_ VGND VGND VPWR VPWR fd._3599_ sky130_fd_sc_hd__xnor2_1
XFILLER_252_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5485_ fd._3917_ fd._0559_ VGND VGND VPWR VPWR fd._0561_ sky130_fd_sc_hd__or2_1
XFILLER_113_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7224_ fd._2468_ fd._2313_ VGND VGND VPWR VPWR fd._2473_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4436_ fd._1913_ fd._3529_ fd._3200_ VGND VGND VPWR VPWR fd._3530_ sky130_fd_sc_hd__mux2_1
XFILLER_113_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7155_ fd._2389_ fd._2393_ fd._2394_ fd._2395_ fd._2396_ VGND VGND VPWR VPWR fd._2398_
+ sky130_fd_sc_hd__o2111a_1
XFILLER_113_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4367_ fd._3211_ VGND VGND VPWR VPWR fd._3222_ sky130_fd_sc_hd__clkbuf_4
XFILLER_208_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6106_ fd._1104_ fd._1243_ VGND VGND VPWR VPWR fd._1244_ sky130_fd_sc_hd__xnor2_1
XFILLER_35_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_263_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7086_ fd._2250_ fd._2321_ VGND VGND VPWR VPWR fd._2322_ sky130_fd_sc_hd__nand2_4
Xfd._4298_ fd.b\[14\] fd._2452_ VGND VGND VPWR VPWR fd._2463_ sky130_fd_sc_hd__nand2_1
XFILLER_39_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_263_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6037_ fd._1059_ fd._1074_ fd._1167_ VGND VGND VPWR VPWR fd._1168_ sky130_fd_sc_hd__or3_1
XFILLER_50_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7988_ fd._3140_ fd._3180_ VGND VGND VPWR VPWR fd._3314_ sky130_fd_sc_hd__nor2_1
XFILLER_33_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6939_ fd._1975_ fd._1981_ VGND VGND VPWR VPWR fd._2160_ sky130_fd_sc_hd__nand2_1
XFILLER_276_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_274_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_274_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_270_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_249_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_265_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_1545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_281_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_281_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_268_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_267_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5270_ fd._3675_ fd._0323_ VGND VGND VPWR VPWR fd._0324_ sky130_fd_sc_hd__xnor2_1
XTAP_5573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4221_ fd.b\[11\] fd._1561_ VGND VGND VPWR VPWR fd._1616_ sky130_fd_sc_hd__or2_1
XTAP_4861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_251_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4152_ fd.b\[10\] VGND VGND VPWR VPWR fd._0857_ sky130_fd_sc_hd__buf_6
XFILLER_263_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_264_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_223_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_225_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4083_ fd.b\[17\] VGND VGND VPWR VPWR fd._0098_ sky130_fd_sc_hd__inv_2
XFILLER_229_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_264_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_225_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7911_ fd._1507_ fd._3226_ VGND VGND VPWR VPWR fd._3229_ sky130_fd_sc_hd__nor2_1
XFILLER_149_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._7842_ fd._2951_ VGND VGND VPWR VPWR fd._3153_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_160_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_258_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4985_ fd._3813_ fd._3927_ VGND VGND VPWR VPWR fd._0011_ sky130_fd_sc_hd__or2_1
Xfd._7773_ fd._3076_ VGND VGND VPWR VPWR fd._3077_ sky130_fd_sc_hd__buf_6
XFILLER_118_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6724_ fd._1728_ fd._1922_ fd._1917_ VGND VGND VPWR VPWR fd._1923_ sky130_fd_sc_hd__mux2_1
XFILLER_144_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_275_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6655_ fd._1431_ fd._1846_ VGND VGND VPWR VPWR fd._1848_ sky130_fd_sc_hd__or2_1
XFILLER_144_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_271_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5606_ fd._0500_ fd._0693_ fd._0614_ VGND VGND VPWR VPWR fd._0694_ sky130_fd_sc_hd__mux2_1
XFILLER_119_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6586_ fd._1397_ fd._1769_ fd._1771_ fd._1585_ VGND VGND VPWR VPWR fd._1772_ sky130_fd_sc_hd__a211o_1
XFILLER_99_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_263_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5537_ fd._0443_ fd._0445_ VGND VGND VPWR VPWR fd._0618_ sky130_fd_sc_hd__and2_1
XFILLER_80_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8256_ net75 net8 VGND VGND VPWR VPWR fd.b\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_269_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5468_ fd._0347_ VGND VGND VPWR VPWR fd._0542_ sky130_fd_sc_hd__clkinv_2
XFILLER_41_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_255_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4419_ fd._0252_ fd._3512_ VGND VGND VPWR VPWR fd._3513_ sky130_fd_sc_hd__nand2_1
XFILLER_187_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7207_ fd._2284_ fd._2286_ VGND VGND VPWR VPWR fd._2455_ sky130_fd_sc_hd__nor2_1
XFILLER_132_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._8187_ net74 fd.mc\[11\] VGND VGND VPWR VPWR fd.c\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_54_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5399_ fd._0456_ fd._0411_ VGND VGND VPWR VPWR fd._0466_ sky130_fd_sc_hd__nand2_1
XFILLER_255_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7138_ fd._2250_ fd._2321_ fd._2378_ fd._2369_ VGND VGND VPWR VPWR fd._2379_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_54_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_282_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_281_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_1663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_1614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_282_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7069_ fd._1632_ fd._2301_ VGND VGND VPWR VPWR fd._2303_ sky130_fd_sc_hd__nor2_1
XFILLER_23_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_274_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1044 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_project_wrapper_103 VGND VGND VPWR VPWR user_project_wrapper_103/HI io_oeb[25]
+ sky130_fd_sc_hd__conb_1
XFILLER_259_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4770_ fd.b\[3\] fd._3686_ VGND VGND VPWR VPWR fd._3864_ sky130_fd_sc_hd__or2_1
Xuser_project_wrapper_114 VGND VGND VPWR VPWR user_project_wrapper_114/HI io_oeb[36]
+ sky130_fd_sc_hd__conb_1
XFILLER_86_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_125 VGND VGND VPWR VPWR user_project_wrapper_125/HI la_data_out[3]
+ sky130_fd_sc_hd__conb_1
XFILLER_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_272_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_project_wrapper_136 VGND VGND VPWR VPWR user_project_wrapper_136/HI la_data_out[14]
+ sky130_fd_sc_hd__conb_1
XFILLER_56_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_project_wrapper_147 VGND VGND VPWR VPWR user_project_wrapper_147/HI la_data_out[25]
+ sky130_fd_sc_hd__conb_1
XFILLER_181_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_158 VGND VGND VPWR VPWR user_project_wrapper_158/HI la_data_out[36]
+ sky130_fd_sc_hd__conb_1
XFILLER_177_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_project_wrapper_169 VGND VGND VPWR VPWR user_project_wrapper_169/HI la_data_out[47]
+ sky130_fd_sc_hd__conb_1
XFILLER_29_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6440_ fd._1609_ fd._1610_ VGND VGND VPWR VPWR fd._1611_ sky130_fd_sc_hd__nor2_1
XFILLER_269_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_268_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_1576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6371_ fd._1534_ VGND VGND VPWR VPWR fd._1535_ sky130_fd_sc_hd__clkinvlp_2
XTAP_6060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_284_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8110_ fd.b\[23\] fd.a\[23\] VGND VGND VPWR VPWR fd._3425_ sky130_fd_sc_hd__and2b_1
XFILLER_231_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._5322_ fd._0288_ fd._0380_ VGND VGND VPWR VPWR fd._0381_ sky130_fd_sc_hd__nand2_1
XFILLER_27_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_271_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._8041_ fd._3370_ fd._3371_ VGND VGND VPWR VPWR fd._3372_ sky130_fd_sc_hd__nor2_1
XFILLER_114_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5253_ fd._0105_ fd._0134_ VGND VGND VPWR VPWR fd._0305_ sky130_fd_sc_hd__and2_1
XFILLER_36_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4204_ fd._0780_ fd._1418_ fd._1220_ VGND VGND VPWR VPWR fd._1429_ sky130_fd_sc_hd__mux2_1
XFILLER_266_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5184_ fd._0036_ fd._0055_ VGND VGND VPWR VPWR fd._0229_ sky130_fd_sc_hd__xor2_1
XFILLER_52_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_263_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4135_ fd.a\[15\] fd.b\[15\] VGND VGND VPWR VPWR fd._0670_ sky130_fd_sc_hd__or2b_1
XFILLER_166_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_1601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._7825_ fd._3132_ fd._3133_ VGND VGND VPWR VPWR fd._3135_ sky130_fd_sc_hd__and2b_1
XFILLER_277_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7756_ fd._3026_ fd._3034_ fd._3055_ fd._3058_ VGND VGND VPWR VPWR fd._3059_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_69_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4968_ fd._3828_ fd._3921_ VGND VGND VPWR VPWR fd._4064_ sky130_fd_sc_hd__nor2_1
XFILLER_195_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6707_ fd._1852_ fd._1900_ fd._1904_ VGND VGND VPWR VPWR fd._1905_ sky130_fd_sc_hd__a21o_1
XFILLER_160_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4899_ fd._3883_ fd._3992_ VGND VGND VPWR VPWR fd._3993_ sky130_fd_sc_hd__and2_1
Xfd._7687_ fd._2790_ fd._2982_ fd._2875_ VGND VGND VPWR VPWR fd._2983_ sky130_fd_sc_hd__mux2_1
XFILLER_275_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6638_ fd._1632_ fd._1828_ VGND VGND VPWR VPWR fd._1829_ sky130_fd_sc_hd__nand2_1
XFILLER_173_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6569_ fd._1582_ fd._1592_ VGND VGND VPWR VPWR fd._1753_ sky130_fd_sc_hd__and2b_1
XFILLER_143_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._8239_ net69 net25 VGND VGND VPWR VPWR fd.a\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_278_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_250_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_1595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5940_ fd._0867_ fd._1060_ fd._1047_ VGND VGND VPWR VPWR fd._1061_ sky130_fd_sc_hd__mux2_1
XFILLER_187_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5871_ fd._0858_ fd._0874_ fd._0984_ VGND VGND VPWR VPWR fd._0985_ sky130_fd_sc_hd__and3_2
XFILLER_179_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7610_ fd._2709_ fd._2897_ fd._2875_ VGND VGND VPWR VPWR fd._2898_ sky130_fd_sc_hd__mux2_1
Xfd._4822_ fd._3908_ fd._3913_ fd._3915_ VGND VGND VPWR VPWR fd._3916_ sky130_fd_sc_hd__a21o_1
XFILLER_31_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4753_ fd._3846_ VGND VGND VPWR VPWR fd._3847_ sky130_fd_sc_hd__inv_2
XFILLER_157_1638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7541_ fd._2680_ fd._2821_ fd._2818_ VGND VGND VPWR VPWR fd._2822_ sky130_fd_sc_hd__a21oi_1
XFILLER_5_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4684_ fd.b\[21\] fd._3776_ VGND VGND VPWR VPWR fd._3778_ sky130_fd_sc_hd__or2_1
Xfd._7472_ fd._2552_ fd._2745_ VGND VGND VPWR VPWR fd._2746_ sky130_fd_sc_hd__nand2_1
XFILLER_29_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_272_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6423_ fd._1015_ fd._1581_ VGND VGND VPWR VPWR fd._1592_ sky130_fd_sc_hd__or2_1
XFILLER_284_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._6354_ fd._1335_ fd._1514_ fd._1515_ fd._1165_ VGND VGND VPWR VPWR fd._1516_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_68_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_256_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5305_ fd._3833_ fd._0166_ VGND VGND VPWR VPWR fd._0363_ sky130_fd_sc_hd__xnor2_1
Xfd._6285_ fd._1293_ fd._1289_ VGND VGND VPWR VPWR fd._1441_ sky130_fd_sc_hd__and2b_1
XFILLER_133_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5236_ fd._0187_ fd._0286_ fd._0269_ VGND VGND VPWR VPWR fd._0287_ sky130_fd_sc_hd__mux2_1
XFILLER_209_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8024_ fd._2076_ fd._3337_ fd._3350_ fd._1666_ VGND VGND VPWR VPWR fd._3353_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_92_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5167_ fd._0200_ fd._0206_ fd._0209_ fd._0210_ VGND VGND VPWR VPWR fd._0211_ sky130_fd_sc_hd__a211o_1
XFILLER_224_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4118_ fd.a\[6\] VGND VGND VPWR VPWR fd._0483_ sky130_fd_sc_hd__inv_2
XFILLER_244_1644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_225_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_269_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5098_ fd._0113_ fd._0119_ fd._0132_ fd._0133_ fd._0134_ VGND VGND VPWR VPWR fd._0135_
+ sky130_fd_sc_hd__o311ai_2
XFILLER_189_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_1675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7808_ fd._1661_ fd._3115_ VGND VGND VPWR VPWR fd._3116_ sky130_fd_sc_hd__and2_1
XFILLER_10_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7739_ fd._2849_ fd._2830_ VGND VGND VPWR VPWR fd._3040_ sky130_fd_sc_hd__nor2_1
XFILLER_279_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_249_1500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_221_ fd.c\[13\] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_1
XFILLER_180_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_1504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_8710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_256_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_8743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_254_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_266_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_250_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6070_ fd._1199_ fd._1203_ fd._1169_ VGND VGND VPWR VPWR fd._1204_ sky130_fd_sc_hd__mux2_1
XFILLER_74_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_262_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5021_ fd._0046_ fd._0039_ fd._0049_ VGND VGND VPWR VPWR fd._0050_ sky130_fd_sc_hd__o21ba_1
XTAP_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_261_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1615 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6972_ fd._1930_ VGND VGND VPWR VPWR fd._2196_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_186_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5923_ fd._0862_ fd._1041_ fd._0861_ VGND VGND VPWR VPWR fd._1042_ sky130_fd_sc_hd__o21ai_2
XFILLER_119_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5854_ fd._0965_ fd._0889_ VGND VGND VPWR VPWR fd._0966_ sky130_fd_sc_hd__nand2_1
XFILLER_255_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4805_ fd._3888_ fd._3893_ fd._3894_ fd._3895_ fd._3898_ VGND VGND VPWR VPWR fd._3899_
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_143_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._5785_ fd._0000_ fd._0889_ VGND VGND VPWR VPWR fd._0891_ sky130_fd_sc_hd__or2_1
XFILLER_142_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7524_ fd._2703_ fd._2801_ fd._2802_ VGND VGND VPWR VPWR fd._2803_ sky130_fd_sc_hd__a21o_1
Xfd._4736_ fd._3726_ fd._3787_ VGND VGND VPWR VPWR fd._3830_ sky130_fd_sc_hd__nand2_1
XFILLER_233_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_269_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7455_ fd._2718_ fd._2725_ fd._2726_ VGND VGND VPWR VPWR fd._2728_ sky130_fd_sc_hd__a21oi_1
Xfd._4667_ fd._3600_ fd._3619_ fd._3604_ VGND VGND VPWR VPWR fd._3761_ sky130_fd_sc_hd__o21a_1
XFILLER_233_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6406_ fd._0427_ fd._1571_ VGND VGND VPWR VPWR fd._1574_ sky130_fd_sc_hd__nand2_1
XFILLER_170_1657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_284_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_256_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4598_ fd._3689_ fd._3691_ fd._3538_ VGND VGND VPWR VPWR fd._3692_ sky130_fd_sc_hd__a21o_1
XFILLER_229_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7386_ fd._1286_ fd._2651_ VGND VGND VPWR VPWR fd._2652_ sky130_fd_sc_hd__or2_1
XFILLER_9_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_1670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6337_ fd._1434_ fd._1497_ VGND VGND VPWR VPWR fd._1498_ sky130_fd_sc_hd__nand2_1
XFILLER_151_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6268_ fd._1349_ VGND VGND VPWR VPWR fd._1422_ sky130_fd_sc_hd__buf_6
XFILLER_77_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8007_ fd._3334_ fd._3198_ fd._3116_ VGND VGND VPWR VPWR fd._3335_ sky130_fd_sc_hd__o21ba_1
XFILLER_240_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5219_ fd._0242_ fd._0244_ VGND VGND VPWR VPWR fd._0268_ sky130_fd_sc_hd__nand2_2
XFILLER_38_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6199_ fd._1327_ fd._1334_ VGND VGND VPWR VPWR fd._1346_ sky130_fd_sc_hd__nor2_1
XFILLER_129_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_279_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_251_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_255_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_261_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_262_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5570_ fd._0553_ VGND VGND VPWR VPWR fd._0654_ sky130_fd_sc_hd__clkinv_2
XFILLER_124_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4521_ fd._2804_ fd._3145_ VGND VGND VPWR VPWR fd._3615_ sky130_fd_sc_hd__or2b_1
XTAP_7872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_1643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4452_ fd._3497_ fd._3490_ VGND VGND VPWR VPWR fd._3546_ sky130_fd_sc_hd__or2b_1
Xfd._7240_ fd._2301_ fd._2490_ fd._2423_ VGND VGND VPWR VPWR fd._2491_ sky130_fd_sc_hd__mux2_1
XFILLER_6_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4383_ fd._2199_ fd._2276_ fd._3387_ fd._2265_ VGND VGND VPWR VPWR fd._3397_ sky130_fd_sc_hd__o31a_1
XFILLER_238_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7171_ fd._2123_ fd._2414_ fd._2323_ VGND VGND VPWR VPWR fd._2415_ sky130_fd_sc_hd__mux2_1
XFILLER_254_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6122_ fd._0916_ fd._1260_ VGND VGND VPWR VPWR fd._1261_ sky130_fd_sc_hd__or2_1
XFILLER_81_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6053_ fd._1184_ VGND VGND VPWR VPWR fd._1185_ sky130_fd_sc_hd__inv_2
XFILLER_222_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_262_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5004_ fd._3802_ fd._0030_ fd._3961_ VGND VGND VPWR VPWR fd._0031_ sky130_fd_sc_hd__mux2_1
XFILLER_59_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_222_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_1636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6955_ fd._2063_ fd._2108_ fd._2109_ fd._2110_ fd._2112_ VGND VGND VPWR VPWR fd._2178_
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_198_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5906_ fd._0995_ fd._0996_ fd._0997_ fd._1023_ VGND VGND VPWR VPWR fd._1024_ sky130_fd_sc_hd__o31a_1
XFILLER_175_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6886_ fd._2083_ fd._2095_ fd._2099_ fd._2101_ VGND VGND VPWR VPWR fd._2102_ sky130_fd_sc_hd__o31a_1
XFILLER_200_1344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5837_ fd._0716_ fd._0902_ VGND VGND VPWR VPWR fd._0948_ sky130_fd_sc_hd__nand2_1
XFILLER_128_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5768_ fd._0871_ fd._0856_ VGND VGND VPWR VPWR fd._0872_ sky130_fd_sc_hd__nand2_1
XFILLER_103_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7507_ fd._2784_ VGND VGND VPWR VPWR fd._2785_ sky130_fd_sc_hd__clkinvlp_2
Xfd._4719_ fd._1253_ fd._3812_ VGND VGND VPWR VPWR fd._3813_ sky130_fd_sc_hd__and2_1
XFILLER_142_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5699_ fd._0775_ fd._0795_ fd._0794_ VGND VGND VPWR VPWR fd._0796_ sky130_fd_sc_hd__and3_1
XFILLER_130_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_269_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7438_ fd._2585_ fd._2677_ fd._2708_ VGND VGND VPWR VPWR fd._2709_ sky130_fd_sc_hd__a21oi_1
XFILLER_131_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_272_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7369_ fd._2434_ fd._2464_ fd._2631_ VGND VGND VPWR VPWR fd._2633_ sky130_fd_sc_hd__a21oi_1
XFILLER_29_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_272_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_281_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_279_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_282_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_251_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6740_ fd._0504_ fd._1940_ VGND VGND VPWR VPWR fd._1941_ sky130_fd_sc_hd__or2_1
XFILLER_157_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_258_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_9060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._6671_ fd._1661_ fd._1648_ fd._1658_ VGND VGND VPWR VPWR fd._1865_ sky130_fd_sc_hd__or3_1
XFILLER_176_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5622_ fd._0490_ fd._0710_ fd._0614_ VGND VGND VPWR VPWR fd._0711_ sky130_fd_sc_hd__mux2_1
XFILLER_171_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5553_ fd._0465_ fd._0481_ fd._0612_ fd._0634_ VGND VGND VPWR VPWR fd._0635_ sky130_fd_sc_hd__a31o_1
XFILLER_124_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4504_ fd._2903_ fd._3597_ fd._3222_ VGND VGND VPWR VPWR fd._3598_ sky130_fd_sc_hd__mux2_1
XFILLER_230_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5484_ fd._0291_ fd._0558_ fd._0452_ VGND VGND VPWR VPWR fd._0559_ sky130_fd_sc_hd__mux2_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7223_ fd._2244_ fd._2471_ fd._2423_ VGND VGND VPWR VPWR fd._2472_ sky130_fd_sc_hd__mux2_1
XFILLER_152_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4435_ fd._3527_ fd._3528_ VGND VGND VPWR VPWR fd._3529_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_254_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_269_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4366_ fd._3200_ VGND VGND VPWR VPWR fd._3211_ sky130_fd_sc_hd__buf_6
Xfd._7154_ fd._1722_ fd._2344_ VGND VGND VPWR VPWR fd._2396_ sky130_fd_sc_hd__xnor2_1
XFILLER_66_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6105_ fd._1111_ fd._1109_ VGND VGND VPWR VPWR fd._1243_ sky130_fd_sc_hd__nor2_1
XFILLER_187_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4297_ fd._0736_ fd._2441_ fd._1220_ VGND VGND VPWR VPWR fd._2452_ sky130_fd_sc_hd__mux2_1
XFILLER_223_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7085_ fd._2297_ fd._2314_ fd._2317_ fd._2319_ VGND VGND VPWR VPWR fd._2321_ sky130_fd_sc_hd__o31a_2
XFILLER_35_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6036_ fd._1079_ fd._1072_ fd._1162_ fd._1166_ VGND VGND VPWR VPWR fd._1167_ sky130_fd_sc_hd__and4b_1
XFILLER_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_277_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7987_ fd._3309_ fd._3312_ fd._3239_ VGND VGND VPWR VPWR fd._3313_ sky130_fd_sc_hd__mux2_1
XFILLER_206_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6938_ fd._1965_ VGND VGND VPWR VPWR fd._2159_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_135_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6869_ fd._2076_ fd._2082_ VGND VGND VPWR VPWR fd._2083_ sky130_fd_sc_hd__nor2_1
XFILLER_151_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_274_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_274_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_252_1573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_281_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_281_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_253_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_268_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_267_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_267_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_276_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4220_ fd._0538_ fd._1594_ fd._1220_ VGND VGND VPWR VPWR fd._1605_ sky130_fd_sc_hd__mux2_1
XFILLER_188_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4151_ fd.b\[11\] VGND VGND VPWR VPWR fd._0846_ sky130_fd_sc_hd__clkinv_4
XFILLER_236_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_1531 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_264_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_251_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4082_ fd._0076_ fd.a\[18\] VGND VGND VPWR VPWR fd._0087_ sky130_fd_sc_hd__nor2_1
XFILLER_205_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7910_ fd._2863_ fd._3220_ VGND VGND VPWR VPWR fd._3228_ sky130_fd_sc_hd__nor2_1
XFILLER_231_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_1540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._7841_ fd._2533_ fd._3151_ VGND VGND VPWR VPWR fd._3152_ sky130_fd_sc_hd__and2_1
XFILLER_125_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7772_ fd._3075_ VGND VGND VPWR VPWR fd._3076_ sky130_fd_sc_hd__buf_6
XFILLER_121_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4984_ fd._3817_ fd._3926_ VGND VGND VPWR VPWR fd._0009_ sky130_fd_sc_hd__nand2_1
XFILLER_157_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6723_ fd._1920_ fd._1921_ VGND VGND VPWR VPWR fd._1922_ sky130_fd_sc_hd__or2_1
XFILLER_201_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1 fd._3405_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_258_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6654_ fd._1843_ fd._1845_ fd._1720_ VGND VGND VPWR VPWR fd._1846_ sky130_fd_sc_hd__mux2_1
XFILLER_132_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_259_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5605_ fd._0690_ fd._0691_ VGND VGND VPWR VPWR fd._0693_ sky130_fd_sc_hd__nand2_1
XFILLER_141_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6585_ fd._0437_ fd._1626_ fd._1644_ fd._1718_ VGND VGND VPWR VPWR fd._1771_ sky130_fd_sc_hd__and4_1
XFILLER_112_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5536_ fd._0616_ VGND VGND VPWR VPWR fd._0617_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_132_1500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8255_ net71 net7 VGND VGND VPWR VPWR fd.b\[15\] sky130_fd_sc_hd__dfxtp_2
XFILLER_239_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5467_ fd._3716_ VGND VGND VPWR VPWR fd._0541_ sky130_fd_sc_hd__buf_6
XFILLER_67_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7206_ fd._2439_ fd._2453_ fd._1494_ VGND VGND VPWR VPWR fd._2454_ sky130_fd_sc_hd__a21o_1
XFILLER_82_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4418_ fd._1825_ fd._3511_ fd._3200_ VGND VGND VPWR VPWR fd._3512_ sky130_fd_sc_hd__mux2_1
XFILLER_27_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8186_ net76 fd.mc\[10\] VGND VGND VPWR VPWR fd.c\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5398_ fd._0455_ fd._0460_ fd._0464_ VGND VGND VPWR VPWR fd._0465_ sky130_fd_sc_hd__o21a_1
XFILLER_187_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_1620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7137_ fd._2377_ fd._2186_ VGND VGND VPWR VPWR fd._2378_ sky130_fd_sc_hd__and2_1
XFILLER_148_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4349_ fd._2573_ fd._2661_ fd._2716_ fd._3002_ fd._3013_ VGND VGND VPWR VPWR fd._3024_
+ sky130_fd_sc_hd__o41a_1
XFILLER_208_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_282_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._7068_ fd._1632_ fd._2301_ VGND VGND VPWR VPWR fd._2302_ sky130_fd_sc_hd__and2_1
XFILLER_39_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6019_ fd._0965_ fd._1140_ fd._1147_ VGND VGND VPWR VPWR fd._1148_ sky130_fd_sc_hd__mux2_1
XFILLER_22_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_276_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_274_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_249_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_259_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_104 VGND VGND VPWR VPWR user_project_wrapper_104/HI io_oeb[26]
+ sky130_fd_sc_hd__conb_1
XFILLER_115_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_115 VGND VGND VPWR VPWR user_project_wrapper_115/HI io_oeb[37]
+ sky130_fd_sc_hd__conb_1
Xuser_project_wrapper_126 VGND VGND VPWR VPWR user_project_wrapper_126/HI la_data_out[4]
+ sky130_fd_sc_hd__conb_1
XFILLER_86_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_137 VGND VGND VPWR VPWR user_project_wrapper_137/HI la_data_out[15]
+ sky130_fd_sc_hd__conb_1
XFILLER_31_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_project_wrapper_148 VGND VGND VPWR VPWR user_project_wrapper_148/HI la_data_out[26]
+ sky130_fd_sc_hd__conb_1
XFILLER_253_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_159 VGND VGND VPWR VPWR user_project_wrapper_159/HI la_data_out[37]
+ sky130_fd_sc_hd__conb_1
XFILLER_257_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_253_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput60 net60 VGND VGND VPWR VPWR io_out[4] sky130_fd_sc_hd__buf_2
XFILLER_116_1517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6370_ fd._1351_ fd._1419_ fd._1533_ VGND VGND VPWR VPWR fd._1534_ sky130_fd_sc_hd__mux2_1
XTAP_6050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5321_ fd._0000_ fd._0287_ VGND VGND VPWR VPWR fd._0380_ sky130_fd_sc_hd__nand2_1
XTAP_6083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_284_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._8040_ fd._3208_ fd._3093_ VGND VGND VPWR VPWR fd._3371_ sky130_fd_sc_hd__and2b_1
XFILLER_23_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5252_ fd._0113_ fd._0119_ fd._0132_ fd._0133_ VGND VGND VPWR VPWR fd._0304_ sky130_fd_sc_hd__o31a_1
XTAP_5393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_270_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4203_ fd._0813_ fd._1407_ VGND VGND VPWR VPWR fd._1418_ sky130_fd_sc_hd__xnor2_1
XFILLER_263_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5183_ fd._0070_ fd._0211_ fd._0226_ fd._0227_ VGND VGND VPWR VPWR fd._0228_ sky130_fd_sc_hd__a31o_1
XFILLER_184_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4134_ fd.b\[15\] fd.a\[15\] VGND VGND VPWR VPWR fd._0659_ sky130_fd_sc_hd__and2b_1
XFILLER_264_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_260_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_264_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_260_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7824_ fd._1722_ fd._3131_ VGND VGND VPWR VPWR fd._3133_ sky130_fd_sc_hd__nand2_1
XFILLER_191_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7755_ fd._2863_ fd._3023_ fd._3056_ VGND VGND VPWR VPWR fd._3058_ sky130_fd_sc_hd__a21o_1
Xfd._4967_ fd._3832_ fd._3920_ VGND VGND VPWR VPWR fd._4063_ sky130_fd_sc_hd__nand2_1
XFILLER_118_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6706_ fd._1903_ VGND VGND VPWR VPWR fd._1904_ sky130_fd_sc_hd__clkinv_4
XFILLER_195_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7686_ fd._2978_ fd._2981_ VGND VGND VPWR VPWR fd._2982_ sky130_fd_sc_hd__xnor2_1
XFILLER_12_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4898_ fd._3867_ fd._3991_ fd._3959_ VGND VGND VPWR VPWR fd._3992_ sky130_fd_sc_hd__mux2_1
XFILLER_47_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6637_ fd._1714_ fd._1827_ fd._1813_ VGND VGND VPWR VPWR fd._1828_ sky130_fd_sc_hd__mux2_1
XFILLER_173_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_1644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6568_ fd._1589_ fd._1591_ VGND VGND VPWR VPWR fd._1752_ sky130_fd_sc_hd__nor2_1
XFILLER_141_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5519_ fd._0594_ fd._0597_ VGND VGND VPWR VPWR fd._0598_ sky130_fd_sc_hd__xnor2_1
XFILLER_41_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6499_ fd._1675_ fd._1481_ VGND VGND VPWR VPWR fd._1676_ sky130_fd_sc_hd__xnor2_1
XFILLER_45_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_214_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._8238_ net68 net24 VGND VGND VPWR VPWR fd.a\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_41_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8169_ fd._3473_ fd._3482_ VGND VGND VPWR VPWR fd._3484_ sky130_fd_sc_hd__or2_1
XFILLER_15_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_270_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_282_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_242_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_266_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5870_ fd._0886_ fd._0979_ fd._0983_ fd._0873_ VGND VGND VPWR VPWR fd._0984_ sky130_fd_sc_hd__o211ai_2
XFILLER_173_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4821_ fd._0846_ fd._3914_ VGND VGND VPWR VPWR fd._3915_ sky130_fd_sc_hd__nor2_1
XFILLER_139_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7540_ fd._2682_ fd._2820_ VGND VGND VPWR VPWR fd._2821_ sky130_fd_sc_hd__nand2_1
Xfd._4752_ fd._3469_ fd._3845_ VGND VGND VPWR VPWR fd._3846_ sky130_fd_sc_hd__nor2_1
XFILLER_155_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_1519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_269_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7471_ fd._0318_ fd._2550_ VGND VGND VPWR VPWR fd._2745_ sky130_fd_sc_hd__nand2_1
XFILLER_138_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4683_ fd._3773_ fd._3776_ VGND VGND VPWR VPWR fd._3777_ sky130_fd_sc_hd__and2_1
XFILLER_155_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6422_ fd._1397_ fd._1588_ fd._1590_ VGND VGND VPWR VPWR fd._1591_ sky130_fd_sc_hd__o21a_1
XFILLER_269_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_268_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_284_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6353_ fd._1336_ fd._1514_ VGND VGND VPWR VPWR fd._1515_ sky130_fd_sc_hd__xor2_1
XFILLER_283_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_284_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5304_ fd._0350_ fd._0356_ fd._0358_ fd._0360_ VGND VGND VPWR VPWR fd._0361_ sky130_fd_sc_hd__a211o_1
XFILLER_83_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6284_ fd._1241_ fd._1283_ VGND VGND VPWR VPWR fd._1439_ sky130_fd_sc_hd__nand2_1
XTAP_5190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8023_ fd._1661_ fd._3348_ fd._3351_ VGND VGND VPWR VPWR fd._3352_ sky130_fd_sc_hd__o21ba_1
XFILLER_114_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5235_ fd._0182_ fd._0284_ VGND VGND VPWR VPWR fd._0286_ sky130_fd_sc_hd__xnor2_1
XFILLER_188_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5166_ fd._1352_ fd._0069_ VGND VGND VPWR VPWR fd._0210_ sky130_fd_sc_hd__nor2_1
XFILLER_52_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4117_ fd._0461_ fd._0241_ fd._0263_ VGND VGND VPWR VPWR fd._0472_ sky130_fd_sc_hd__o21ba_1
XFILLER_240_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5097_ fd._3883_ fd._0103_ VGND VGND VPWR VPWR fd._0134_ sky130_fd_sc_hd__or2_1
XFILLER_225_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_269_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_277_1443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7807_ fd._2983_ fd._3114_ fd._3076_ VGND VGND VPWR VPWR fd._3115_ sky130_fd_sc_hd__mux2_1
XFILLER_192_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5999_ fd._1118_ fd._1123_ VGND VGND VPWR VPWR fd._1126_ sky130_fd_sc_hd__nor2_1
XFILLER_195_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7738_ fd._3038_ VGND VGND VPWR VPWR fd._3039_ sky130_fd_sc_hd__inv_2
XFILLER_69_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_279_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7669_ fd._2942_ VGND VGND VPWR VPWR fd._2963_ sky130_fd_sc_hd__inv_2
XFILLER_121_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_249_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_220_ fd.c\[12\] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_1
XFILLER_168_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_8711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5020_ fd._0047_ fd._0048_ fd._3946_ VGND VGND VPWR VPWR fd._0049_ sky130_fd_sc_hd__mux2_1
XFILLER_228_1629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6971_ fd._2152_ fd._2158_ fd._2192_ fd._2193_ fd._2194_ VGND VGND VPWR VPWR fd._2195_
+ sky130_fd_sc_hd__o311a_1
XFILLER_124_1627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5922_ fd._1040_ fd._0981_ fd._0869_ VGND VGND VPWR VPWR fd._1041_ sky130_fd_sc_hd__o21ai_1
XFILLER_204_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5853_ fd._0000_ VGND VGND VPWR VPWR fd._0965_ sky130_fd_sc_hd__buf_6
XFILLER_31_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_1559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4804_ fd._3897_ VGND VGND VPWR VPWR fd._3898_ sky130_fd_sc_hd__inv_2
XFILLER_115_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5784_ fd._0735_ fd._0888_ fd._0848_ VGND VGND VPWR VPWR fd._0889_ sky130_fd_sc_hd__mux2_1
XFILLER_127_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7523_ fd._1645_ fd._2697_ VGND VGND VPWR VPWR fd._2802_ sky130_fd_sc_hd__nor2_1
XFILLER_5_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4735_ fd._3723_ fd._3727_ VGND VGND VPWR VPWR fd._3829_ sky130_fd_sc_hd__xnor2_1
XFILLER_103_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_272_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_272_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._7454_ fd._2566_ fd._2717_ VGND VGND VPWR VPWR fd._2726_ sky130_fd_sc_hd__and2_1
Xfd._4666_ fd._3610_ VGND VGND VPWR VPWR fd._3760_ sky130_fd_sc_hd__clkinv_2
XFILLER_269_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6405_ fd._0427_ fd._1571_ VGND VGND VPWR VPWR fd._1573_ sky130_fd_sc_hd__nor2_1
XFILLER_9_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7385_ fd._2449_ fd._2649_ fd._2506_ VGND VGND VPWR VPWR fd._2651_ sky130_fd_sc_hd__mux2_1
Xfd._4597_ fd._3537_ fd._3222_ VGND VGND VPWR VPWR fd._3691_ sky130_fd_sc_hd__nor2_1
XFILLER_151_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_256_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6336_ fd._0594_ fd._1433_ VGND VGND VPWR VPWR fd._1497_ sky130_fd_sc_hd__or2_1
XFILLER_84_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_284_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_272_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6267_ fd._1303_ fd._1420_ VGND VGND VPWR VPWR fd._1421_ sky130_fd_sc_hd__xnor2_1
XFILLER_37_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8006_ fd._3127_ fd._3197_ VGND VGND VPWR VPWR fd._3334_ sky130_fd_sc_hd__and2_1
XFILLER_52_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5218_ fd._0228_ fd._0234_ VGND VGND VPWR VPWR fd._0267_ sky130_fd_sc_hd__xnor2_1
XFILLER_225_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6198_ fd._1314_ fd._1321_ VGND VGND VPWR VPWR fd._1345_ sky130_fd_sc_hd__or2_1
XFILLER_240_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._5149_ fd._4069_ fd._4062_ fd._4068_ VGND VGND VPWR VPWR fd._0191_ sky130_fd_sc_hd__and3_1
XFILLER_209_1551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_279_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_279_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1495 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_279_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_1560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_251_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_261_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_1586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_1548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4520_ fd._2793_ VGND VGND VPWR VPWR fd._3614_ sky130_fd_sc_hd__clkinv_2
XTAP_7851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_285_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4451_ fd._3510_ fd._3514_ fd._3543_ fd._3544_ fd._3508_ VGND VGND VPWR VPWR fd._3545_
+ sky130_fd_sc_hd__o311a_1
XFILLER_215_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7170_ fd._2228_ fd._2413_ VGND VGND VPWR VPWR fd._2414_ sky130_fd_sc_hd__nor2_1
XFILLER_43_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4382_ fd._2144_ fd._2221_ VGND VGND VPWR VPWR fd._3387_ sky130_fd_sc_hd__nor2_1
XFILLER_266_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6121_ fd._1086_ fd._1259_ fd._1169_ VGND VGND VPWR VPWR fd._1260_ sky130_fd_sc_hd__mux2_1
XFILLER_171_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_267_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_253_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6052_ fd._1178_ fd._1183_ VGND VGND VPWR VPWR fd._1184_ sky130_fd_sc_hd__xnor2_1
XFILLER_165_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_262_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5003_ fd._0027_ fd._0029_ VGND VGND VPWR VPWR fd._0030_ sky130_fd_sc_hd__xor2_1
XFILLER_179_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_1659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6954_ fd._2044_ fd._2047_ VGND VGND VPWR VPWR fd._2176_ sky130_fd_sc_hd__or2_1
XFILLER_119_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5905_ fd._3537_ fd._0829_ VGND VGND VPWR VPWR fd._1023_ sky130_fd_sc_hd__xnor2_1
XFILLER_174_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._6885_ fd._0382_ fd._2098_ VGND VGND VPWR VPWR fd._2101_ sky130_fd_sc_hd__or2_1
XFILLER_50_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5836_ fd._0541_ fd._0946_ VGND VGND VPWR VPWR fd._0947_ sky130_fd_sc_hd__or2_1
XFILLER_200_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5767_ fd._0786_ fd._0855_ VGND VGND VPWR VPWR fd._0871_ sky130_fd_sc_hd__nand2_1
XFILLER_172_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7506_ fd._2725_ fd._2783_ VGND VGND VPWR VPWR fd._2784_ sky130_fd_sc_hd__nand2_1
Xfd._4718_ fd._3745_ fd._3810_ fd._3800_ fd._3811_ VGND VGND VPWR VPWR fd._3812_ sky130_fd_sc_hd__a31oi_2
XFILLER_153_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5698_ fd._0776_ fd._0767_ VGND VGND VPWR VPWR fd._0795_ sky130_fd_sc_hd__nand2_1
XFILLER_9_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7437_ fd._2582_ fd._2670_ fd._2675_ VGND VGND VPWR VPWR fd._2708_ sky130_fd_sc_hd__and3_1
XFILLER_285_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4649_ fd._3645_ fd._3742_ VGND VGND VPWR VPWR fd._3743_ sky130_fd_sc_hd__nand2_1
XFILLER_229_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7368_ fd._2434_ fd._2464_ fd._2631_ VGND VGND VPWR VPWR fd._2632_ sky130_fd_sc_hd__and3_1
XFILLER_69_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_268_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6319_ fd._4055_ fd._1280_ VGND VGND VPWR VPWR fd._1478_ sky130_fd_sc_hd__xnor2_1
XFILLER_211_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_272_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7299_ fd._1970_ fd._2423_ fd._2498_ fd._2504_ fd._2555_ VGND VGND VPWR VPWR fd._2556_
+ sky130_fd_sc_hd__a41o_1
XFILLER_44_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_225_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_285_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_279_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_1592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_257_1688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_1639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6670_ fd._0726_ fd._1863_ VGND VGND VPWR VPWR fd._1864_ sky130_fd_sc_hd__nor2_1
XTAP_9050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5621_ fd._0492_ fd._0709_ VGND VGND VPWR VPWR fd._0710_ sky130_fd_sc_hd__xnor2_1
XFILLER_67_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_258_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5552_ fd._0624_ fd._0633_ VGND VGND VPWR VPWR fd._0634_ sky130_fd_sc_hd__or2b_1
XFILLER_158_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4503_ fd._3596_ fd._2991_ VGND VGND VPWR VPWR fd._3597_ sky130_fd_sc_hd__xnor2_1
XTAP_7681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._8271_ net69 net25 VGND VGND VPWR VPWR fd.b\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_267_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5483_ fd._0361_ fd._0557_ VGND VGND VPWR VPWR fd._0558_ sky130_fd_sc_hd__nand2_1
XFILLER_6_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._7222_ fd._2470_ VGND VGND VPWR VPWR fd._2471_ sky130_fd_sc_hd__clkinv_2
Xfd._4434_ fd._1935_ fd._1990_ VGND VGND VPWR VPWR fd._3528_ sky130_fd_sc_hd__nand2_1
XFILLER_230_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_282_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7153_ fd._2135_ fd._2392_ VGND VGND VPWR VPWR fd._2395_ sky130_fd_sc_hd__or2_1
XFILLER_113_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4365_ fd._3156_ fd._3178_ fd._3189_ VGND VGND VPWR VPWR fd._3200_ sky130_fd_sc_hd__a21o_4
XFILLER_26_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6104_ fd._0726_ fd._1240_ VGND VGND VPWR VPWR fd._1241_ sky130_fd_sc_hd__or2_1
XFILLER_130_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._7084_ fd._2310_ fd._2318_ fd._2317_ VGND VGND VPWR VPWR fd._2319_ sky130_fd_sc_hd__or3_1
XFILLER_39_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4296_ fd._2419_ fd._2430_ VGND VGND VPWR VPWR fd._2441_ sky130_fd_sc_hd__xor2_1
XFILLER_207_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6035_ fd._0482_ fd._1161_ fd._1164_ VGND VGND VPWR VPWR fd._1166_ sky130_fd_sc_hd__o21ai_1
XFILLER_165_1535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7986_ fd._3190_ fd._3311_ VGND VGND VPWR VPWR fd._3312_ sky130_fd_sc_hd__xnor2_1
XFILLER_277_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6937_ fd._1559_ fd._2157_ VGND VGND VPWR VPWR fd._2158_ sky130_fd_sc_hd__and2_1
XFILLER_190_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6868_ fd._2079_ fd._2080_ fd._1969_ fd._2081_ VGND VGND VPWR VPWR fd._2082_ sky130_fd_sc_hd__o31a_1
XFILLER_89_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5819_ fd._3658_ VGND VGND VPWR VPWR fd._0928_ sky130_fd_sc_hd__buf_6
XFILLER_200_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6799_ fd._1795_ fd._1794_ VGND VGND VPWR VPWR fd._2006_ sky130_fd_sc_hd__or2b_1
XFILLER_143_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_273_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_281_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_263_1692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_253_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4150_ fd._0417_ fd._0505_ fd._0648_ fd._0824_ VGND VGND VPWR VPWR fd._0835_ sky130_fd_sc_hd__a211o_1
XTAP_4896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4081_ fd.b\[18\] VGND VGND VPWR VPWR fd._0076_ sky130_fd_sc_hd__inv_2
XFILLER_32_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._7840_ fd._2941_ fd._3150_ fd._3075_ VGND VGND VPWR VPWR fd._3151_ sky130_fd_sc_hd__mux2_1
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7771_ fd._3074_ fd._3038_ fd._3050_ fd._3060_ VGND VGND VPWR VPWR fd._3075_ sky130_fd_sc_hd__a31o_4
XFILLER_258_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4983_ fd._4070_ fd._0006_ fd._0007_ fd._0004_ VGND VGND VPWR VPWR fd._0008_ sky130_fd_sc_hd__a211o_1
XFILLER_199_1664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6722_ fd._1731_ fd._1919_ VGND VGND VPWR VPWR fd._1921_ sky130_fd_sc_hd__nor2_1
XFILLER_157_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_2 fd._3695_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6653_ fd._1690_ fd._1844_ VGND VGND VPWR VPWR fd._1845_ sky130_fd_sc_hd__xnor2_1
XFILLER_126_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5604_ fd._0536_ fd._0689_ VGND VGND VPWR VPWR fd._0691_ sky130_fd_sc_hd__or2_1
XFILLER_154_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_263_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6584_ fd._1626_ fd._1644_ fd._1718_ fd._1768_ VGND VGND VPWR VPWR fd._1769_ sky130_fd_sc_hd__a31o_1
XFILLER_119_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_8190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5535_ fd._0426_ fd._0448_ fd._0614_ VGND VGND VPWR VPWR fd._0616_ sky130_fd_sc_hd__mux2_1
XFILLER_119_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8254_ net71 net6 VGND VGND VPWR VPWR fd.b\[14\] sky130_fd_sc_hd__dfxtp_2
XFILLER_267_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5466_ fd._0492_ fd._0503_ fd._0539_ fd._0489_ VGND VGND VPWR VPWR fd._0540_ sky130_fd_sc_hd__a31oi_2
XFILLER_6_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_255_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_269_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7205_ fd._2447_ fd._2448_ fd._2451_ fd._2444_ VGND VGND VPWR VPWR fd._2453_ sky130_fd_sc_hd__o211ai_2
XFILLER_67_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4417_ fd._1847_ fd._2023_ VGND VGND VPWR VPWR fd._3511_ sky130_fd_sc_hd__xnor2_1
XFILLER_187_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_269_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._8185_ net76 fd.mc\[9\] VGND VGND VPWR VPWR fd.c\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_66_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5397_ fd._0271_ fd._0462_ fd._0463_ VGND VGND VPWR VPWR fd._0464_ sky130_fd_sc_hd__mux2_1
XFILLER_27_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7136_ fd._1585_ VGND VGND VPWR VPWR fd._2377_ sky130_fd_sc_hd__buf_6
XFILLER_270_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4348_ fd._2705_ fd._2639_ fd._3002_ fd._2694_ VGND VGND VPWR VPWR fd._3013_ sky130_fd_sc_hd__a211o_1
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7067_ fd._2053_ fd._2300_ fd._2238_ VGND VGND VPWR VPWR fd._2301_ sky130_fd_sc_hd__mux2_1
Xfd._4279_ fd._2232_ fd._2243_ fd._1220_ VGND VGND VPWR VPWR fd._2254_ sky130_fd_sc_hd__mux2_1
XFILLER_212_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6018_ fd._0965_ fd._1146_ VGND VGND VPWR VPWR fd._1147_ sky130_fd_sc_hd__xnor2_1
XFILLER_282_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7969_ fd._1751_ fd._3286_ fd._3292_ VGND VGND VPWR VPWR fd._3293_ sky130_fd_sc_hd__a21o_1
XFILLER_202_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_249_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_1601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_253_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_1530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_281_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_259_1536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_105 VGND VGND VPWR VPWR user_project_wrapper_105/HI io_oeb[27]
+ sky130_fd_sc_hd__conb_1
XFILLER_177_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_259_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_116 VGND VGND VPWR VPWR user_project_wrapper_116/HI io_out[32]
+ sky130_fd_sc_hd__conb_1
Xuser_project_wrapper_127 VGND VGND VPWR VPWR user_project_wrapper_127/HI la_data_out[5]
+ sky130_fd_sc_hd__conb_1
Xuser_project_wrapper_138 VGND VGND VPWR VPWR user_project_wrapper_138/HI la_data_out[16]
+ sky130_fd_sc_hd__conb_1
XFILLER_108_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_project_wrapper_149 VGND VGND VPWR VPWR user_project_wrapper_149/HI la_data_out[27]
+ sky130_fd_sc_hd__conb_1
XFILLER_194_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput50 net50 VGND VGND VPWR VPWR io_out[24] sky130_fd_sc_hd__buf_2
XFILLER_268_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_1545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput61 net61 VGND VGND VPWR VPWR io_out[5] sky130_fd_sc_hd__buf_2
XFILLER_96_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_268_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_284_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_1580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1591 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5320_ fd._1308_ fd._0378_ VGND VGND VPWR VPWR fd._0379_ sky130_fd_sc_hd__or2_1
XTAP_6073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5251_ fd._0089_ fd._0295_ fd._0302_ VGND VGND VPWR VPWR fd._0303_ sky130_fd_sc_hd__a21o_1
XFILLER_188_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4202_ fd._1396_ fd._0648_ fd._0912_ VGND VGND VPWR VPWR fd._1407_ sky130_fd_sc_hd__o21ai_1
XFILLER_236_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5182_ fd._0224_ fd._0215_ fd._0223_ VGND VGND VPWR VPWR fd._0227_ sky130_fd_sc_hd__o21ba_1
XTAP_4693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4133_ fd._0516_ fd._0560_ fd._0637_ VGND VGND VPWR VPWR fd._0648_ sky130_fd_sc_hd__or3_1
XFILLER_252_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_258_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_1671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7823_ fd._1722_ fd._3131_ VGND VGND VPWR VPWR fd._3132_ sky130_fd_sc_hd__nor2_1
XFILLER_121_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4966_ fd._4054_ fd._3646_ fd._4061_ VGND VGND VPWR VPWR fd._4062_ sky130_fd_sc_hd__mux2_1
Xfd._7754_ fd._2861_ fd._3022_ fd._2877_ VGND VGND VPWR VPWR fd._3056_ sky130_fd_sc_hd__a21o_1
XFILLER_117_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6705_ fd._1848_ fd._1901_ VGND VGND VPWR VPWR fd._1903_ sky130_fd_sc_hd__and2_1
XFILLER_195_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7685_ fd._2979_ fd._2791_ VGND VGND VPWR VPWR fd._2981_ sky130_fd_sc_hd__nor2_1
Xfd._4897_ fd._3868_ fd._3983_ VGND VGND VPWR VPWR fd._3991_ sky130_fd_sc_hd__xnor2_1
XFILLER_86_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6636_ fd._1703_ fd._1826_ VGND VGND VPWR VPWR fd._1827_ sky130_fd_sc_hd__xnor2_1
XFILLER_67_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1607 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._6567_ fd._0427_ VGND VGND VPWR VPWR fd._1751_ sky130_fd_sc_hd__buf_6
XFILLER_119_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5518_ fd._0453_ fd._0596_ VGND VGND VPWR VPWR fd._0597_ sky130_fd_sc_hd__nand2_1
XFILLER_113_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6498_ fd._1470_ fd._1475_ fd._1476_ VGND VGND VPWR VPWR fd._1675_ sky130_fd_sc_hd__o21bai_1
XFILLER_132_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_1686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5449_ fd._0520_ VGND VGND VPWR VPWR fd._0521_ sky130_fd_sc_hd__clkinvlp_2
Xfd._8237_ net68 net22 VGND VGND VPWR VPWR fd.a\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_255_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8168_ fd._3473_ fd._3482_ VGND VGND VPWR VPWR fd._3483_ sky130_fd_sc_hd__nand2_1
XFILLER_23_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7119_ fd._2357_ fd._2349_ VGND VGND VPWR VPWR fd._2358_ sky130_fd_sc_hd__xnor2_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._8099_ fd._0270_ fd._0453_ fd._3411_ VGND VGND VPWR VPWR fd._3419_ sky130_fd_sc_hd__mux2_1
XFILLER_39_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_270_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_282_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1578 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_254_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_266_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_284_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_265_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_281_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4820_ fd._3912_ VGND VGND VPWR VPWR fd._3914_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_122_1566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4751_ fd._3844_ fd._3661_ fd._3787_ VGND VGND VPWR VPWR fd._3845_ sky130_fd_sc_hd__mux2_1
XFILLER_170_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7470_ fd._0821_ fd._2556_ fd._2557_ VGND VGND VPWR VPWR fd._2744_ sky130_fd_sc_hd__a21o_1
XFILLER_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_272_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4682_ fd._3598_ fd._3626_ fd._3774_ fd._3775_ VGND VGND VPWR VPWR fd._3776_ sky130_fd_sc_hd__o22a_1
XFILLER_237_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6421_ fd._3695_ fd._1533_ fd._1211_ VGND VGND VPWR VPWR fd._1590_ sky130_fd_sc_hd__o21ai_2
XFILLER_116_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_268_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6352_ fd._1508_ fd._1329_ fd._1327_ VGND VGND VPWR VPWR fd._1514_ sky130_fd_sc_hd__a21oi_1
XFILLER_81_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5303_ fd._0846_ fd._0359_ VGND VGND VPWR VPWR fd._0360_ sky130_fd_sc_hd__nor2_1
XFILLER_284_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6283_ fd._1294_ fd._1436_ fd._1423_ fd._1437_ VGND VGND VPWR VPWR fd._1438_ sky130_fd_sc_hd__a31o_1
XFILLER_49_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8022_ fd._1666_ fd._3350_ fd._3348_ fd._1661_ VGND VGND VPWR VPWR fd._3351_ sky130_fd_sc_hd__a22o_1
XFILLER_42_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_266_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5234_ fd._0189_ fd._0188_ VGND VGND VPWR VPWR fd._0284_ sky130_fd_sc_hd__or2b_1
XFILLER_237_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5165_ fd._0075_ fd._0199_ fd._0206_ fd._0207_ VGND VGND VPWR VPWR fd._0209_ sky130_fd_sc_hd__o31a_1
XFILLER_184_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_283_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4116_ fd._0450_ fd.a\[4\] VGND VGND VPWR VPWR fd._0461_ sky130_fd_sc_hd__nand2_1
XFILLER_252_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_264_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5096_ fd._3675_ fd._0112_ VGND VGND VPWR VPWR fd._0133_ sky130_fd_sc_hd__or2_1
XFILLER_189_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7806_ fd._2977_ fd._3113_ VGND VGND VPWR VPWR fd._3114_ sky130_fd_sc_hd__xnor2_1
XFILLER_140_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5998_ fd._1124_ VGND VGND VPWR VPWR fd._1125_ sky130_fd_sc_hd__clkinv_4
XFILLER_121_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7737_ fd._3026_ fd._3037_ VGND VGND VPWR VPWR fd._3038_ sky130_fd_sc_hd__nor2_2
Xfd._4949_ fd._3915_ fd._3913_ VGND VGND VPWR VPWR fd._4043_ sky130_fd_sc_hd__and2b_1
XFILLER_160_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7668_ fd._2952_ fd._2957_ fd._2960_ fd._2961_ VGND VGND VPWR VPWR fd._2962_ sky130_fd_sc_hd__o31ai_2
XFILLER_133_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_271_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6619_ fd._1807_ fd._1641_ VGND VGND VPWR VPWR fd._1808_ sky130_fd_sc_hd__and2b_1
XFILLER_271_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7599_ fd._0207_ fd._2884_ VGND VGND VPWR VPWR fd._2886_ sky130_fd_sc_hd__nand2_1
XFILLER_113_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_249_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_250_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_266_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_265_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6970_ fd._2150_ VGND VGND VPWR VPWR fd._2194_ sky130_fd_sc_hd__clkinvlp_2
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5921_ fd._0886_ fd._0979_ VGND VGND VPWR VPWR fd._1040_ sky130_fd_sc_hd__nor2_1
XFILLER_169_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5852_ fd._1308_ fd._0963_ VGND VGND VPWR VPWR fd._0964_ sky130_fd_sc_hd__nor2_1
XFILLER_200_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4803_ fd._3851_ fd._3896_ VGND VGND VPWR VPWR fd._3897_ sky130_fd_sc_hd__nand2_1
XFILLER_155_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5783_ fd._0731_ fd._0887_ VGND VGND VPWR VPWR fd._0888_ sky130_fd_sc_hd__xnor2_1
XFILLER_142_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._4734_ fd._3646_ fd._3827_ VGND VGND VPWR VPWR fd._3828_ sky130_fd_sc_hd__nor2_1
XFILLER_196_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7522_ fd._2707_ fd._2798_ fd._2800_ VGND VGND VPWR VPWR fd._2801_ sky130_fd_sc_hd__a21o_1
XFILLER_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4665_ fd._3757_ fd._3758_ VGND VGND VPWR VPWR fd._3759_ sky130_fd_sc_hd__nand2_1
XFILLER_170_1604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7453_ fd._1173_ fd._2724_ VGND VGND VPWR VPWR fd._2725_ sky130_fd_sc_hd__nand2_1
XFILLER_237_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6404_ fd._1389_ fd._1570_ fd._1533_ VGND VGND VPWR VPWR fd._1571_ sky130_fd_sc_hd__mux2_1
XFILLER_170_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7384_ fd._2647_ fd._2648_ VGND VGND VPWR VPWR fd._2649_ sky130_fd_sc_hd__xor2_1
XFILLER_9_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4596_ fd._3689_ fd._3222_ VGND VGND VPWR VPWR fd._3690_ sky130_fd_sc_hd__nand2_1
XFILLER_190_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6335_ fd._1444_ fd._1493_ fd._1494_ VGND VGND VPWR VPWR fd._1496_ sky130_fd_sc_hd__a21o_1
XFILLER_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._6266_ fd._1338_ fd._1307_ VGND VGND VPWR VPWR fd._1420_ sky130_fd_sc_hd__nor2_1
XFILLER_42_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5217_ fd._0260_ fd._0265_ VGND VGND VPWR VPWR fd._0266_ sky130_fd_sc_hd__xnor2_1
Xfd._8005_ fd._3327_ fd._3330_ fd._3331_ VGND VGND VPWR VPWR fd._3333_ sky130_fd_sc_hd__or3b_1
XFILLER_20_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6197_ fd._1058_ fd._1342_ fd._1048_ VGND VGND VPWR VPWR fd._1344_ sky130_fd_sc_hd__a21boi_1
XFILLER_77_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5148_ fd._0182_ fd._0188_ fd._0189_ VGND VGND VPWR VPWR fd._0190_ sky130_fd_sc_hd__a21oi_1
XFILLER_52_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_283_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._5079_ fd._4006_ fd._4009_ VGND VGND VPWR VPWR fd._0114_ sky130_fd_sc_hd__or2_1
XFILLER_220_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_279_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_261_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_249_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_273_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4450_ fd._0428_ fd._3502_ VGND VGND VPWR VPWR fd._3544_ sky130_fd_sc_hd__or2_1
XFILLER_254_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_1678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_227_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4381_ fd.b\[13\] fd._3365_ VGND VGND VPWR VPWR fd._3376_ sky130_fd_sc_hd__or2_1
XFILLER_281_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_285_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._6120_ fd._1250_ fd._1251_ VGND VGND VPWR VPWR fd._1259_ sky130_fd_sc_hd__xnor2_1
XFILLER_187_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_253_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6051_ fd._1006_ fd._1182_ fd._1169_ VGND VGND VPWR VPWR fd._1183_ sky130_fd_sc_hd__mux2_1
XFILLER_185_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_250_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5002_ fd._0028_ fd._3931_ VGND VGND VPWR VPWR fd._0029_ sky130_fd_sc_hd__nor2_1
XFILLER_206_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6953_ fd._2021_ fd._2026_ fd._2032_ VGND VGND VPWR VPWR fd._2175_ sky130_fd_sc_hd__a21oi_1
XFILLER_148_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5904_ fd._0437_ fd._0849_ VGND VGND VPWR VPWR fd._1021_ sky130_fd_sc_hd__nand2_1
XFILLER_200_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6884_ fd._0382_ fd._2098_ VGND VGND VPWR VPWR fd._2099_ sky130_fd_sc_hd__and2_1
XFILLER_204_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5835_ fd._0705_ fd._0944_ fd._0848_ VGND VGND VPWR VPWR fd._0946_ sky130_fd_sc_hd__mux2_1
XFILLER_174_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_274_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5766_ fd._0863_ fd._0869_ VGND VGND VPWR VPWR fd._0870_ sky130_fd_sc_hd__nand2_1
XFILLER_157_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7505_ fd._1173_ fd._2724_ VGND VGND VPWR VPWR fd._2783_ sky130_fd_sc_hd__or2_1
Xfd._4717_ fd._3644_ fd._3800_ VGND VGND VPWR VPWR fd._3811_ sky130_fd_sc_hd__nor2_1
XFILLER_118_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5697_ fd._0793_ VGND VGND VPWR VPWR fd._0794_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_157_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7436_ fd._1872_ fd._2706_ VGND VGND VPWR VPWR fd._2707_ sky130_fd_sc_hd__or2_1
Xfd._4648_ fd._2584_ fd._3644_ VGND VGND VPWR VPWR fd._3742_ sky130_fd_sc_hd__nand2_1
XFILLER_269_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4579_ fd._3519_ fd._3672_ fd._3624_ VGND VGND VPWR VPWR fd._3673_ sky130_fd_sc_hd__mux2_1
Xfd._7367_ fd._2426_ fd._2466_ VGND VGND VPWR VPWR fd._2631_ sky130_fd_sc_hd__nor2_1
XFILLER_29_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_285_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_284_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_285_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_272_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_268_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6318_ fd._1470_ fd._1475_ fd._1476_ VGND VGND VPWR VPWR fd._1477_ sky130_fd_sc_hd__o21ba_1
XFILLER_84_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7298_ fd._2498_ fd._2504_ fd._2554_ VGND VGND VPWR VPWR fd._2555_ sky130_fd_sc_hd__a21oi_1
XFILLER_272_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._6249_ fd._0318_ fd._1391_ fd._1398_ fd._1400_ VGND VGND VPWR VPWR fd._1401_ sky130_fd_sc_hd__a22o_1
XFILLER_53_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_279_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_1492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_263_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_243_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_262_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_1614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_9062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5620_ fd._0503_ fd._0539_ VGND VGND VPWR VPWR fd._0709_ sky130_fd_sc_hd__nand2_1
XTAP_9084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_259_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5551_ fd._0632_ fd._0444_ VGND VGND VPWR VPWR fd._0633_ sky130_fd_sc_hd__nand2_1
XFILLER_140_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4502_ fd.b\[18\] fd._2947_ fd._3595_ VGND VGND VPWR VPWR fd._3596_ sky130_fd_sc_hd__a21bo_1
XTAP_7682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5482_ fd._0358_ fd._0556_ VGND VGND VPWR VPWR fd._0557_ sky130_fd_sc_hd__nand2_1
Xfd._8270_ net68 net24 VGND VGND VPWR VPWR fd.b\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_285_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_267_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4433_ fd._1979_ fd._3526_ VGND VGND VPWR VPWR fd._3527_ sky130_fd_sc_hd__and2_1
XTAP_6981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7221_ fd._2469_ fd._2316_ VGND VGND VPWR VPWR fd._2470_ sky130_fd_sc_hd__xor2_1
XTAP_6992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_266_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_267_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_254_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4364_ fd._1231_ VGND VGND VPWR VPWR fd._3189_ sky130_fd_sc_hd__clkinv_2
Xfd._7152_ fd._2346_ fd._2339_ VGND VGND VPWR VPWR fd._2394_ sky130_fd_sc_hd__and2b_1
XFILLER_66_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_254_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6103_ fd._1123_ fd._1239_ fd._1223_ VGND VGND VPWR VPWR fd._1240_ sky130_fd_sc_hd__mux2_1
XFILLER_47_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7083_ fd._2312_ fd._2302_ VGND VGND VPWR VPWR fd._2318_ sky130_fd_sc_hd__nor2_1
XFILLER_19_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4295_ fd._0802_ fd._1407_ fd._0791_ VGND VGND VPWR VPWR fd._2430_ sky130_fd_sc_hd__a21oi_1
XFILLER_35_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6034_ fd._0883_ fd._1163_ fd._1047_ VGND VGND VPWR VPWR fd._1164_ sky130_fd_sc_hd__mux2_1
XFILLER_165_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_223_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._7985_ fd._3196_ fd._3195_ VGND VGND VPWR VPWR fd._3311_ sky130_fd_sc_hd__or2b_1
XFILLER_147_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6936_ fd._2153_ fd._2156_ fd._2115_ VGND VGND VPWR VPWR fd._2157_ sky130_fd_sc_hd__mux2_1
XFILLER_276_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6867_ fd._1868_ fd._1969_ VGND VGND VPWR VPWR fd._2081_ sky130_fd_sc_hd__nand2_1
XFILLER_50_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5818_ fd._0926_ VGND VGND VPWR VPWR fd._0927_ sky130_fd_sc_hd__clkinv_4
XFILLER_11_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6798_ fd._1933_ fd._1997_ fd._2003_ fd._2004_ VGND VGND VPWR VPWR fd._2005_ sky130_fd_sc_hd__a31o_1
XFILLER_89_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5749_ fd._0755_ fd._0756_ fd._0763_ fd._0779_ VGND VGND VPWR VPWR fd._0851_ sky130_fd_sc_hd__a31o_1
XFILLER_137_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._7419_ fd._2055_ fd._2687_ VGND VGND VPWR VPWR fd._2688_ sky130_fd_sc_hd__nor2_1
XFILLER_69_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_257_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_279_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_279_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4080_ fd._0032_ fd._0054_ VGND VGND VPWR VPWR fd._0065_ sky130_fd_sc_hd__nor2_1
XFILLER_205_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7770_ fd._0131_ fd._3073_ fd._3020_ VGND VGND VPWR VPWR fd._3074_ sky130_fd_sc_hd__mux2_1
XFILLER_61_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4982_ fd._1253_ fd._3971_ VGND VGND VPWR VPWR fd._0007_ sky130_fd_sc_hd__nor2_1
XFILLER_12_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_258_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_1507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6721_ fd._1731_ fd._1919_ VGND VGND VPWR VPWR fd._1920_ sky130_fd_sc_hd__and2_1
XFILLER_195_1518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_3 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._6652_ fd._1698_ fd._1697_ VGND VGND VPWR VPWR fd._1844_ sky130_fd_sc_hd__or2b_1
XFILLER_6_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5603_ fd._0536_ fd._0689_ VGND VGND VPWR VPWR fd._0690_ sky130_fd_sc_hd__nand2_1
XFILLER_158_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._6583_ fd._1590_ fd._1765_ VGND VGND VPWR VPWR fd._1768_ sky130_fd_sc_hd__nand2_1
XFILLER_4_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5534_ fd._0613_ VGND VGND VPWR VPWR fd._0614_ sky130_fd_sc_hd__buf_6
XFILLER_154_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._8253_ net71 net5 VGND VGND VPWR VPWR fd.b\[13\] sky130_fd_sc_hd__dfxtp_2
XFILLER_112_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5465_ fd._0525_ fd._0531_ fd._0532_ fd._0534_ fd._0537_ VGND VGND VPWR VPWR fd._0539_
+ sky130_fd_sc_hd__a2111o_1
XFILLER_227_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7204_ fd._2450_ VGND VGND VPWR VPWR fd._2451_ sky130_fd_sc_hd__clkinvlp_2
Xfd._4416_ fd._3508_ fd._3509_ VGND VGND VPWR VPWR fd._3510_ sky130_fd_sc_hd__nand2_1
Xfd._5396_ fd._0279_ fd._0449_ fd._0277_ VGND VGND VPWR VPWR fd._0463_ sky130_fd_sc_hd__o21ai_1
Xfd._8184_ net76 fd.mc\[8\] VGND VGND VPWR VPWR fd.c\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4347_ fd._2980_ fd._2991_ VGND VGND VPWR VPWR fd._3002_ sky130_fd_sc_hd__or2_1
XFILLER_255_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7135_ fd._1764_ fd._2179_ fd._2250_ fd._2321_ VGND VGND VPWR VPWR fd._2376_ sky130_fd_sc_hd__o211a_1
XFILLER_187_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4278_ fd._1385_ fd._0626_ VGND VGND VPWR VPWR fd._2243_ sky130_fd_sc_hd__xnor2_1
Xuser_project_wrapper_90 VGND VGND VPWR VPWR user_project_wrapper_90/HI io_oeb[12]
+ sky130_fd_sc_hd__conb_1
Xfd._7066_ fd._2299_ fd._2106_ VGND VGND VPWR VPWR fd._2300_ sky130_fd_sc_hd__xnor2_1
XFILLER_39_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6017_ fd._1141_ fd._1145_ fd._1046_ VGND VGND VPWR VPWR fd._1146_ sky130_fd_sc_hd__mux2_1
XFILLER_247_1699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7968_ fd._2533_ fd._3291_ VGND VGND VPWR VPWR fd._3292_ sky130_fd_sc_hd__and2_1
XFILLER_124_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_276_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6919_ fd._1943_ fd._2137_ VGND VGND VPWR VPWR fd._2138_ sky130_fd_sc_hd__xnor2_1
XFILLER_136_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7899_ fd._3048_ fd._3049_ VGND VGND VPWR VPWR fd._3216_ sky130_fd_sc_hd__and2_1
XFILLER_11_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_274_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_253_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_265_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_246_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1580 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_1608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_259_1548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_106 VGND VGND VPWR VPWR user_project_wrapper_106/HI io_oeb[28]
+ sky130_fd_sc_hd__conb_1
XFILLER_154_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_117 VGND VGND VPWR VPWR user_project_wrapper_117/HI io_out[33]
+ sky130_fd_sc_hd__conb_1
XFILLER_147_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_project_wrapper_128 VGND VGND VPWR VPWR user_project_wrapper_128/HI la_data_out[6]
+ sky130_fd_sc_hd__conb_1
XFILLER_68_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_139 VGND VGND VPWR VPWR user_project_wrapper_139/HI la_data_out[17]
+ sky130_fd_sc_hd__conb_1
XFILLER_29_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput40 net40 VGND VGND VPWR VPWR io_out[15] sky130_fd_sc_hd__buf_2
XFILLER_190_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput51 net51 VGND VGND VPWR VPWR io_out[25] sky130_fd_sc_hd__buf_2
XFILLER_29_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput62 net62 VGND VGND VPWR VPWR io_out[6] sky130_fd_sc_hd__buf_2
XTAP_6030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_253_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_1412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5250_ fd._0089_ fd._0295_ fd._0301_ VGND VGND VPWR VPWR fd._0302_ sky130_fd_sc_hd__o21a_1
XTAP_5373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4201_ fd._1385_ VGND VGND VPWR VPWR fd._1396_ sky130_fd_sc_hd__inv_2
XTAP_4661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5181_ fd._0218_ fd._0225_ VGND VGND VPWR VPWR fd._0226_ sky130_fd_sc_hd__and2_1
XFILLER_188_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4132_ fd._0593_ fd._0626_ VGND VGND VPWR VPWR fd._0637_ sky130_fd_sc_hd__nand2_1
XTAP_3971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_260_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_242_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7822_ fd._2970_ fd._3130_ fd._3075_ VGND VGND VPWR VPWR fd._3131_ sky130_fd_sc_hd__mux2_1
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_1558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_277_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7753_ fd._2856_ fd._3054_ VGND VGND VPWR VPWR fd._3055_ sky130_fd_sc_hd__xor2_1
XFILLER_9_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4965_ fd._4055_ fd._4059_ VGND VGND VPWR VPWR fd._4061_ sky130_fd_sc_hd__xnor2_1
XFILLER_195_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6704_ fd._1431_ fd._1846_ VGND VGND VPWR VPWR fd._1901_ sky130_fd_sc_hd__nand2_1
XFILLER_274_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7684_ fd._2326_ fd._2790_ VGND VGND VPWR VPWR fd._2979_ sky130_fd_sc_hd__nor2_1
Xfd._4896_ fd._3988_ fd._3989_ VGND VGND VPWR VPWR fd._3990_ sky130_fd_sc_hd__nand2_1
XFILLER_12_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6635_ fd._1716_ fd._1709_ VGND VGND VPWR VPWR fd._1826_ sky130_fd_sc_hd__or2_1
XFILLER_126_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6566_ fd._1559_ fd._1749_ VGND VGND VPWR VPWR fd._1750_ sky130_fd_sc_hd__and2_1
XFILLER_134_1619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_271_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_253_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_1632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5517_ fd._1264_ fd._0595_ VGND VGND VPWR VPWR fd._0596_ sky130_fd_sc_hd__xnor2_1
XFILLER_80_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_268_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6497_ fd._1645_ fd._1668_ fd._1673_ VGND VGND VPWR VPWR fd._1674_ sky130_fd_sc_hd__mux2_1
XFILLER_234_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8236_ net68 net21 VGND VGND VPWR VPWR fd.a\[28\] sky130_fd_sc_hd__dfxtp_1
Xfd._5448_ fd._0312_ fd._0519_ VGND VGND VPWR VPWR fd._0520_ sky130_fd_sc_hd__nor2_1
XFILLER_28_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_255_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8167_ fd._3478_ fd._3481_ VGND VGND VPWR VPWR fd._3482_ sky130_fd_sc_hd__xnor2_1
XFILLER_82_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5379_ fd._3695_ fd._0425_ VGND VGND VPWR VPWR fd._0444_ sky130_fd_sc_hd__nor2_1
XFILLER_167_1417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_255_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_270_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7118_ fd._2190_ fd._2348_ VGND VGND VPWR VPWR fd._2357_ sky130_fd_sc_hd__and2_1
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8098_ fd._3418_ VGND VGND VPWR VPWR fd.mc\[16\] sky130_fd_sc_hd__clkbuf_1
XFILLER_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_282_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7049_ fd._2280_ fd._2099_ VGND VGND VPWR VPWR fd._2281_ sky130_fd_sc_hd__nor2_1
XFILLER_54_1609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_254_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_278_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_219_1554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_274_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_265_1596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1670 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_1578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4750_ fd._3710_ fd._3843_ VGND VGND VPWR VPWR fd._3844_ sky130_fd_sc_hd__nand2_1
XFILLER_196_1668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4681_ fd._3600_ fd._3623_ VGND VGND VPWR VPWR fd._3775_ sky130_fd_sc_hd__or2b_1
XFILLER_177_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6420_ fd._1397_ fd._1588_ VGND VGND VPWR VPWR fd._1589_ sky130_fd_sc_hd__and2_1
XFILLER_155_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6351_ fd._1505_ fd._1511_ fd._1512_ VGND VGND VPWR VPWR fd._1513_ sky130_fd_sc_hd__a21o_1
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_268_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5302_ fd._0355_ VGND VGND VPWR VPWR fd._0359_ sky130_fd_sc_hd__inv_2
XFILLER_110_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6282_ fd._1236_ fd._1422_ VGND VGND VPWR VPWR fd._1437_ sky130_fd_sc_hd__nor2_1
XTAP_5170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_260_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._8021_ fd._3115_ fd._3349_ fd._3239_ VGND VGND VPWR VPWR fd._3350_ sky130_fd_sc_hd__mux2_1
XFILLER_252_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5233_ fd._1264_ fd._0282_ VGND VGND VPWR VPWR fd._0283_ sky130_fd_sc_hd__or2_1
XFILLER_188_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_251_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5164_ fd._0076_ VGND VGND VPWR VPWR fd._0207_ sky130_fd_sc_hd__buf_8
XFILLER_252_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4115_ fd._0219_ VGND VGND VPWR VPWR fd._0450_ sky130_fd_sc_hd__clkinv_8
XFILLER_205_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._5095_ fd._3869_ fd._0118_ fd._0126_ fd._0130_ VGND VGND VPWR VPWR fd._0132_ sky130_fd_sc_hd__o211a_1
XFILLER_33_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_277_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7805_ fd._2987_ fd._2984_ VGND VGND VPWR VPWR fd._3113_ sky130_fd_sc_hd__and2b_1
XFILLER_118_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5997_ fd._1118_ fd._1123_ VGND VGND VPWR VPWR fd._1124_ sky130_fd_sc_hd__nand2_1
XFILLER_195_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7736_ fd._3034_ fd._3036_ VGND VGND VPWR VPWR fd._3037_ sky130_fd_sc_hd__nand2_1
XFILLER_121_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._4948_ fd._4035_ fd._4039_ fd._4041_ VGND VGND VPWR VPWR fd._4042_ sky130_fd_sc_hd__a21o_1
XFILLER_133_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7667_ fd._2751_ fd._2951_ VGND VGND VPWR VPWR fd._2961_ sky130_fd_sc_hd__or2_1
XFILLER_47_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4879_ fd._3888_ fd._3893_ fd._3895_ VGND VGND VPWR VPWR fd._3973_ sky130_fd_sc_hd__o21ai_1
XFILLER_218_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6618_ fd._1631_ fd._1806_ fd._1643_ VGND VGND VPWR VPWR fd._1807_ sky130_fd_sc_hd__a21o_1
XFILLER_173_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._7598_ fd._0207_ fd._2884_ VGND VGND VPWR VPWR fd._2885_ sky130_fd_sc_hd__or2_1
XFILLER_59_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6549_ fd._1729_ fd._1730_ VGND VGND VPWR VPWR fd._1731_ sky130_fd_sc_hd__nor2_1
XFILLER_214_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8219_ net73 net3 VGND VGND VPWR VPWR fd.a\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_255_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_271_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_282_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_260_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_259_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_266_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_265_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_267_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_1636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_1601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_261_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_261_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_261_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5920_ fd._1035_ fd._1038_ VGND VGND VPWR VPWR fd._1039_ sky130_fd_sc_hd__xnor2_1
XFILLER_187_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5851_ fd._0961_ fd._0962_ fd._0848_ VGND VGND VPWR VPWR fd._0963_ sky130_fd_sc_hd__mux2_1
XFILLER_161_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4802_ fd._2155_ fd._3850_ VGND VGND VPWR VPWR fd._3896_ sky130_fd_sc_hd__nand2_1
XFILLER_31_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5782_ fd._0738_ fd._0737_ VGND VGND VPWR VPWR fd._0887_ sky130_fd_sc_hd__or2b_1
XFILLER_115_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_259_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7521_ fd._2703_ fd._2799_ VGND VGND VPWR VPWR fd._2800_ sky130_fd_sc_hd__nand2_1
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4733_ fd._3825_ fd._3788_ fd._3826_ VGND VGND VPWR VPWR fd._3827_ sky130_fd_sc_hd__o21ai_1
XFILLER_154_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7452_ fd._2719_ fd._2723_ fd._2676_ VGND VGND VPWR VPWR fd._2724_ sky130_fd_sc_hd__mux2_1
Xfd._4664_ fd._3628_ fd._3752_ fd._3756_ VGND VGND VPWR VPWR fd._3758_ sky130_fd_sc_hd__nand3_1
XFILLER_269_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6403_ fd._1567_ fd._1569_ VGND VGND VPWR VPWR fd._1570_ sky130_fd_sc_hd__xnor2_1
XFILLER_25_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_284_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7383_ fd._2439_ fd._2451_ VGND VGND VPWR VPWR fd._2648_ sky130_fd_sc_hd__nand2_1
XFILLER_96_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_269_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4595_ fd.b\[0\] VGND VGND VPWR VPWR fd._3689_ sky130_fd_sc_hd__buf_6
XFILLER_57_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_284_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_250_1662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfd._6334_ fd._0098_ VGND VGND VPWR VPWR fd._1494_ sky130_fd_sc_hd__buf_6
XFILLER_81_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_284_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6265_ fd._1414_ fd._1417_ VGND VGND VPWR VPWR fd._1419_ sky130_fd_sc_hd__xnor2_1
XFILLER_49_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8004_ fd._1173_ fd._3326_ fd._3329_ fd._2566_ VGND VGND VPWR VPWR fd._3331_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_246_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._5216_ fd._0261_ fd._0264_ VGND VGND VPWR VPWR fd._0265_ sky130_fd_sc_hd__and2b_1
XFILLER_253_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6196_ fd._1048_ fd._1342_ VGND VGND VPWR VPWR fd._1343_ sky130_fd_sc_hd__and2b_1
XFILLER_65_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_252_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5147_ fd._1297_ fd._0187_ VGND VGND VPWR VPWR fd._0189_ sky130_fd_sc_hd__and2_1
XFILLER_224_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5078_ fd._3675_ fd._0112_ VGND VGND VPWR VPWR fd._0113_ sky130_fd_sc_hd__xnor2_2
XFILLER_33_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_277_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7719_ fd._3009_ fd._3015_ fd._3016_ fd._3017_ VGND VGND VPWR VPWR fd._3018_ sky130_fd_sc_hd__o211a_1
XFILLER_279_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_255_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_263_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_284_1224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_278_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1662 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_1337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_254_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_285_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_266_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4380_ fd._1506_ fd._3211_ fd._3354_ VGND VGND VPWR VPWR fd._3365_ sky130_fd_sc_hd__o21ai_1
XFILLER_215_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_266_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_253_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_281_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._6050_ fd._1180_ fd._1181_ VGND VGND VPWR VPWR fd._1182_ sky130_fd_sc_hd__xnor2_1
XFILLER_111_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5001_ fd._3803_ VGND VGND VPWR VPWR fd._0028_ sky130_fd_sc_hd__inv_2
XFILLER_267_1499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_261_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._6952_ fd._1958_ fd._2173_ VGND VGND VPWR VPWR fd._2174_ sky130_fd_sc_hd__and2_1
XFILLER_124_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfd._5903_ fd._1015_ fd._1019_ VGND VGND VPWR VPWR fd._1020_ sky130_fd_sc_hd__nand2_1
XFILLER_147_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._6883_ fd._1887_ fd._2097_ fd._1917_ VGND VGND VPWR VPWR fd._2098_ sky130_fd_sc_hd__mux2_1
XFILLER_50_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5834_ fd._0700_ fd._0943_ VGND VGND VPWR VPWR fd._0944_ sky130_fd_sc_hd__xnor2_1
XFILLER_162_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5765_ fd._0768_ fd._0867_ VGND VGND VPWR VPWR fd._0869_ sky130_fd_sc_hd__or2_1
XFILLER_171_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7504_ fd._2780_ VGND VGND VPWR VPWR fd._2781_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_282_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._4716_ fd._3743_ fd._3809_ VGND VGND VPWR VPWR fd._3810_ sky130_fd_sc_hd__nand2_1
XFILLER_48_1541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5696_ fd._0785_ fd._0792_ VGND VGND VPWR VPWR fd._0793_ sky130_fd_sc_hd__or2_1
XFILLER_174_1560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_276_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_269_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7435_ fd._2590_ fd._2704_ fd._2677_ VGND VGND VPWR VPWR fd._2706_ sky130_fd_sc_hd__mux2_1
Xfd._4647_ fd._1297_ fd._3740_ VGND VGND VPWR VPWR fd._3741_ sky130_fd_sc_hd__or2_1
XFILLER_9_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._7366_ fd._2627_ VGND VGND VPWR VPWR fd._2630_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_9_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4578_ fd._3522_ fd._3541_ VGND VGND VPWR VPWR fd._3672_ sky130_fd_sc_hd__xnor2_1
XFILLER_97_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6317_ fd._1118_ fd._1474_ VGND VGND VPWR VPWR fd._1476_ sky130_fd_sc_hd__and2_1
XFILLER_238_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._7297_ fd._2381_ fd._2553_ VGND VGND VPWR VPWR fd._2554_ sky130_fd_sc_hd__nand2_1
XFILLER_84_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6248_ fd._1397_ fd._1393_ fd._1395_ fd._0632_ fd._1399_ VGND VGND VPWR VPWR fd._1400_
+ sky130_fd_sc_hd__o32ai_1
XFILLER_168_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6179_ fd._1304_ fd._1161_ VGND VGND VPWR VPWR fd._1324_ sky130_fd_sc_hd__or2_1
XFILLER_225_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_279_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_257_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_251_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_279_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_1625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_263_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_250_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_1522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_9074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_9085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_8373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5550_ fd._4011_ VGND VGND VPWR VPWR fd._0632_ sky130_fd_sc_hd__buf_4
XTAP_8384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4501_ fd.b\[18\] fd._2947_ fd._3585_ VGND VGND VPWR VPWR fd._3595_ sky130_fd_sc_hd__o21bai_1
XTAP_7661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._5481_ fd._0350_ fd._0356_ fd._0360_ VGND VGND VPWR VPWR fd._0556_ sky130_fd_sc_hd__a21o_1
XFILLER_79_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._7220_ fd._2312_ fd._2468_ fd._2308_ VGND VGND VPWR VPWR fd._2469_ sky130_fd_sc_hd__o21a_1
XFILLER_94_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4432_ fd.b\[0\] fd._3525_ VGND VGND VPWR VPWR fd._3526_ sky130_fd_sc_hd__or2_1
XFILLER_6_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7151_ fd._2135_ fd._2392_ VGND VGND VPWR VPWR fd._2393_ sky130_fd_sc_hd__and2_1
Xfd._4363_ fd._3167_ fd._1198_ fd._1187_ VGND VGND VPWR VPWR fd._3178_ sky130_fd_sc_hd__mux2_1
XFILLER_43_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6102_ fd._1117_ fd._1238_ VGND VGND VPWR VPWR fd._1239_ sky130_fd_sc_hd__xnor2_1
XFILLER_81_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7082_ fd._2239_ fd._2316_ VGND VGND VPWR VPWR fd._2317_ sky130_fd_sc_hd__nand2_1
Xfd._4294_ fd._0747_ fd._0769_ VGND VGND VPWR VPWR fd._2419_ sky130_fd_sc_hd__nor2_1
XFILLER_228_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6033_ fd._1064_ fd._0975_ VGND VGND VPWR VPWR fd._1163_ sky130_fd_sc_hd__xor2_1
XFILLER_262_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_280_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7984_ fd._3194_ VGND VGND VPWR VPWR fd._3309_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_206_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6935_ fd._2154_ fd._2145_ VGND VGND VPWR VPWR fd._2156_ sky130_fd_sc_hd__xnor2_1
XFILLER_198_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6866_ fd._1879_ fd._1884_ fd._2077_ VGND VGND VPWR VPWR fd._2080_ sky130_fd_sc_hd__and3_1
XFILLER_147_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5817_ fd._0917_ fd._0915_ VGND VGND VPWR VPWR fd._0926_ sky130_fd_sc_hd__or2b_1
XFILLER_190_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6797_ fd._0343_ fd._2002_ VGND VGND VPWR VPWR fd._2004_ sky130_fd_sc_hd__nor2_1
XFILLER_157_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5748_ fd._0788_ fd._0847_ fd._0849_ VGND VGND VPWR VPWR fd._0850_ sky130_fd_sc_hd__mux2_1
XFILLER_171_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_277_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_256_1690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5679_ fd._0475_ fd._0773_ fd._0651_ VGND VGND VPWR VPWR fd._0774_ sky130_fd_sc_hd__mux2_1
XFILLER_276_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7418_ fd._2508_ fd._2686_ fd._2677_ VGND VGND VPWR VPWR fd._2687_ sky130_fd_sc_hd__mux2_1
XFILLER_285_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_285_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_268_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7349_ fd._2415_ fd._2577_ VGND VGND VPWR VPWR fd._2611_ sky130_fd_sc_hd__nand2_1
XFILLER_84_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_285_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_272_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_285_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_279_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_275_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_279_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_267_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_257_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_257_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_1610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_283_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_270_1665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_249_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_282_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_268_1572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_251_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_264_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4981_ fd._0004_ fd._0005_ VGND VGND VPWR VPWR fd._0006_ sky130_fd_sc_hd__nor2_1
XFILLER_223_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6720_ fd._1736_ fd._1778_ VGND VGND VPWR VPWR fd._1919_ sky130_fd_sc_hd__nor2_1
XFILLER_185_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_258_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_4 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfd._6651_ fd._1696_ VGND VGND VPWR VPWR fd._1843_ sky130_fd_sc_hd__clkinv_2
XFILLER_67_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._5602_ fd._0525_ fd._0531_ fd._0534_ VGND VGND VPWR VPWR fd._0689_ sky130_fd_sc_hd__a21oi_1
XFILLER_271_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfd._6582_ fd._1719_ fd._1763_ fd._1766_ fd._0821_ VGND VGND VPWR VPWR fd._1767_ sky130_fd_sc_hd__o211ai_2
XFILLER_154_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_271_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_8170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_259_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_8192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._5533_ fd._0465_ fd._0481_ fd._0612_ VGND VGND VPWR VPWR fd._0613_ sky130_fd_sc_hd__nand3_2
XFILLER_193_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8252_ net73 net4 VGND VGND VPWR VPWR fd.b\[12\] sky130_fd_sc_hd__dfxtp_2
XFILLER_234_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5464_ fd._0536_ VGND VGND VPWR VPWR fd._0537_ sky130_fd_sc_hd__inv_2
XFILLER_171_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_269_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_267_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7203_ fd._2055_ fd._2449_ VGND VGND VPWR VPWR fd._2450_ sky130_fd_sc_hd__nor2_1
XFILLER_94_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_254_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4415_ fd.b\[6\] fd._3507_ VGND VGND VPWR VPWR fd._3509_ sky130_fd_sc_hd__nand2_1
XFILLER_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._8183_ net77 fd.mc\[7\] VGND VGND VPWR VPWR fd.c\[7\] sky130_fd_sc_hd__dfxtp_1
Xfd._5395_ fd._0271_ fd._0424_ VGND VGND VPWR VPWR fd._0462_ sky130_fd_sc_hd__nand2_1
XFILLER_27_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_282_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_254_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7134_ fd._1958_ fd._2373_ VGND VGND VPWR VPWR fd._2374_ sky130_fd_sc_hd__nand2_1
XFILLER_48_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._4346_ fd._2925_ fd._2958_ VGND VGND VPWR VPWR fd._2991_ sky130_fd_sc_hd__or2b_1
XFILLER_82_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_270_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7065_ fd._1431_ fd._2292_ fd._2107_ VGND VGND VPWR VPWR fd._2299_ sky130_fd_sc_hd__mux2_1
XFILLER_19_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4277_ fd.a\[8\] VGND VGND VPWR VPWR fd._2232_ sky130_fd_sc_hd__clkinv_2
XFILLER_208_1607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_80 VGND VGND VPWR VPWR user_project_wrapper_80/HI io_oeb[2]
+ sky130_fd_sc_hd__conb_1
Xuser_project_wrapper_91 VGND VGND VPWR VPWR user_project_wrapper_91/HI io_oeb[13]
+ sky130_fd_sc_hd__conb_1
XFILLER_34_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfd._6016_ fd._0960_ fd._1144_ VGND VGND VPWR VPWR fd._1145_ sky130_fd_sc_hd__xnor2_1
XFILLER_165_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7967_ fd._3287_ fd._3290_ fd._3239_ VGND VGND VPWR VPWR fd._3291_ sky130_fd_sc_hd__mux2_1
XFILLER_163_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._6918_ fd._1949_ fd._1985_ VGND VGND VPWR VPWR fd._2137_ sky130_fd_sc_hd__nor2_1
XFILLER_135_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_276_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._7898_ fd._3069_ fd._3214_ VGND VGND VPWR VPWR fd._3215_ sky130_fd_sc_hd__xor2_1
XFILLER_15_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6849_ fd._1853_ fd._2060_ fd._2020_ VGND VGND VPWR VPWR fd._2061_ sky130_fd_sc_hd__mux2_1
XFILLER_135_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_254_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_278_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_281_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_1549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_107 VGND VGND VPWR VPWR user_project_wrapper_107/HI io_oeb[29]
+ sky130_fd_sc_hd__conb_1
XFILLER_182_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_project_wrapper_118 VGND VGND VPWR VPWR user_project_wrapper_118/HI io_out[34]
+ sky130_fd_sc_hd__conb_1
XFILLER_154_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xuser_project_wrapper_129 VGND VGND VPWR VPWR user_project_wrapper_129/HI la_data_out[7]
+ sky130_fd_sc_hd__conb_1
XFILLER_68_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_1577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput41 net41 VGND VGND VPWR VPWR io_out[16] sky130_fd_sc_hd__buf_2
XFILLER_123_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput52 net52 VGND VGND VPWR VPWR io_out[26] sky130_fd_sc_hd__buf_2
XFILLER_122_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput63 net63 VGND VGND VPWR VPWR io_out[7] sky130_fd_sc_hd__buf_2
XFILLER_1_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4200_ fd._0417_ fd._0505_ VGND VGND VPWR VPWR fd._1385_ sky130_fd_sc_hd__nand2_1
XFILLER_236_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_252_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5180_ fd._0223_ fd._0224_ VGND VGND VPWR VPWR fd._0225_ sky130_fd_sc_hd__nor2_1
XTAP_4673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_1485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfd._4131_ fd._0604_ fd._0615_ VGND VGND VPWR VPWR fd._0626_ sky130_fd_sc_hd__nor2_1
XFILLER_252_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_260_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7821_ fd._2965_ fd._3129_ VGND VGND VPWR VPWR fd._3130_ sky130_fd_sc_hd__xor2_1
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_277_1605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfd._7752_ fd._3053_ fd._2865_ fd._2864_ VGND VGND VPWR VPWR fd._3054_ sky130_fd_sc_hd__a21o_1
XFILLER_117_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4964_ fd._3920_ fd._4057_ fd._3960_ fd._4058_ VGND VGND VPWR VPWR fd._4059_ sky130_fd_sc_hd__a31o_1
XFILLER_160_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_277_1649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_258_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6703_ fd._1275_ fd._1853_ fd._1898_ fd._0965_ fd._1899_ VGND VGND VPWR VPWR fd._1900_
+ sky130_fd_sc_hd__a221o_1
XFILLER_117_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._7683_ fd._2728_ fd._2786_ VGND VGND VPWR VPWR fd._2978_ sky130_fd_sc_hd__nor2_1
XFILLER_12_1565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._4895_ fd._3669_ fd._3987_ VGND VGND VPWR VPWR fd._3989_ sky130_fd_sc_hd__nand2_1
XFILLER_173_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_275_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6634_ fd._1165_ fd._1823_ VGND VGND VPWR VPWR fd._1824_ sky130_fd_sc_hd__nand2_1
XFILLER_114_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_1677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfd._6565_ fd._1571_ fd._1747_ fd._1719_ VGND VGND VPWR VPWR fd._1749_ sky130_fd_sc_hd__mux2_1
XFILLER_154_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._5516_ fd._0288_ fd._0386_ VGND VGND VPWR VPWR fd._0595_ sky130_fd_sc_hd__nand2_1
XFILLER_98_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfd._6496_ fd._4055_ fd._1672_ VGND VGND VPWR VPWR fd._1673_ sky130_fd_sc_hd__xnor2_1
.ends

